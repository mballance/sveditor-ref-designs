
`include "uvm_macros.svh"

package my_xt_agent_pkg;
	import uvm_pkg::*;
	
	`include "my_xt_config.svh"
	`include "my_xt_seq_item.svh"
	`include "my_xt_driver.svh"
	`include "my_xt_monitor.svh"
	`include "my_xt_seq_base.svh"
	`include "my_xt_agent.svh"
endpackage




// ========== Copyright Header Begin ==========================================
// 
// OpenSPARC T2 Processor File: forcePORstate.vh
// Copyright (C) 1995-2007 Sun Microsystems, Inc. All Rights Reserved
// 4150 Network Circle, Santa Clara, California 95054, U.S.A.
//
// * DO NOT ALTER OR REMOVE COPYRIGHT NOTICES OR THIS FILE HEADER. 
//
// This program is free software; you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation; version 2 of the License.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA
// 
// For the avoidance of doubt, and except that if any non-GPL license 
// choice is available it will apply instead, Sun elects to use only 
// the General Public License version 2 (GPLv2) at this time for any 
// software where a choice of GPL license versions is made 
// available with the language indicating that GPLv2 or any later version 
// may be used, or where a choice of which version of the GPL is applied is 
// otherwise unspecified. 
//
// Please contact Sun Microsystems, Inc., 4150 Network Circle, Santa Clara, 
// CA 95054 USA or visit www.sun.com if you need additional information or 
// have any questions. 
// 
// ========== Copyright Header End ============================================
force tb_top.cpu.ccx.clk_ccx.xcluster_header_left.alatch.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_left.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_left.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_left.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_left.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_left.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_left.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_left.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_left.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.alatch.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.ccx.clk_ccx.xcluster_header_right.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ccx.clk_ccx.xcluster_header_right.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_0.d0_0 value=1111111111111111111111111111111111111111111111111111111111111111 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_0.d0_0.d = 64'b0000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_1.d0_0 value=1111111111111111111111111111111111111111111111111111111111111111 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_1.d0_0.d = 64'b0000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_2.d0_0 value=111111111 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_2.d0_0.d = 9'b000000000;

// instance=tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_3.d0_0 value=111111111 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_3.d0_0.d = 9'b000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl0.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl0.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl1.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl1.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl2.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl2.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl3.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl3.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl4.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl4.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl5.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl5.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl6.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl6.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbl7.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbl7.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr0.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr0.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr1.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr1.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr2.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr2.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr3.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr3.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr4.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr4.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr5.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr5.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr6.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr6.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.cpx.cpx_arbr7.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.cpx.cpx_arbr7.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.bfd0.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd0.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd0.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd0.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd0.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd0.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd0.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd0.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd1.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd1.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd1.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd1.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd1.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd1.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd1.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd1.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd2.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd2.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd2.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd2.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd2.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd2.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd2.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd2.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd3.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd3.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd3.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd3.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd3.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd3.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd3.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd3.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd4.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd4.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd4.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd4.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd4.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd4.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd4.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd4.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd5.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd5.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd5.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd5.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd5.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd5.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd5.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd5.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd6.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd6.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd6.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd6.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd6.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd6.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd6.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd6.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd7.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd7.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd7.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd7.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd7.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd7.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd7.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd7.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_0.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_0.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_1.d0_0 value=1100000000000000000000000000000000000000000000000000000000000011 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_1.d0_0.d = 64'b0011111111111111111111111111111111111111111111111111111111111100;

// instance=tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_2.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_2.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_3.d0_0 value=100000 out=q_l in=d model=msffiz_dp 
force tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_3.d0_0.d = 6'b011111;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl0.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl0.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl1.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl1.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl2.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl2.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl3.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl3.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl4.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl4.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl5.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl5.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl6.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl6.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl7.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl7.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbl8.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbl8.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr0.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr0.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr1.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr1.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr2.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr2.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr3.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr3.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr4.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr4.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr5.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr5.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr6.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr6.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr7.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr7.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.dff_inreg_select.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.dff_inreg_select.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q0.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q0.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q1.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q1.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q2.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q2.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q3.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q3.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q4.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q4.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q5.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q5.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q6.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q6.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q7.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q7.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q8.dff_qfullbar_a.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q8.dff_qfullbar_a.d0_0.d = 1'b1;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.ard.i_dff_qual_atomic_d1.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.ard.i_dff_qual_atomic_d1.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.ccx.pcx.pcx_arbr8.ard.i_dff_req_a.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.ccx.pcx.pcx_arbr8.ard.i_dff_req_a.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.dbg0.db0_clk_header_iol2clk.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.dbg0.db0_clk_header_iol2clk.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.dbg0.rtc.ff_io_sync_en.d0_0 value=10001000110000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.dbg0.rtc.ff_io_sync_en.d0_0.d = 50'b10001000110000000000000000000000000000000000000000;

// instance=tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.dbg1.db1_clk_header_iol2clk.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.dbg1.db1_clk_header_iol2clk.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.dbg1.dbg1_dbgprt.ff_cmp_io_sync_en.d0_0 value=0100010001111000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.dbg1.dbg1_dbgprt.ff_cmp_io_sync_en.d0_0.d = 37'b0100010001111000000000000000000000000;

// instance=tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_0.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_0.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_1.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_1.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_2.d0_0 value=1111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_2.d0_0.d = 22'b1111111111111111111111;

// instance=tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_seq_gen.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_seq_gen.d0_0.d = 2'b11;

// instance=tb_top.cpu.efu.efu_ioclk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.efu.efu_ioclk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.efu.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.efu.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.efu.niu_interface.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.efu.niu_interface.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.efu.niu_interface.ff_mcu_fclrz.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.efu.niu_interface.ff_mcu_fclrz.d0_0.d = 1'b1;

// instance=tb_top.cpu.efu.niu_interface.ff_niu_fclrz.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.efu.niu_interface.ff_niu_fclrz.d0_0.d = 1'b1;

// instance=tb_top.cpu.efu.niu_interface.ff_psr_fclrz.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.efu.niu_interface.ff_psr_fclrz.d0_0.d = 1'b1;

// instance=tb_top.cpu.efu.u_efa_stdc.enable_efa_por_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.efu.u_efa_stdc.enable_efa_por_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b0.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b0.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b0.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b0.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b0.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b0.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b0.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b0.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b0.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b0.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b0.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b0.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b0.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b0.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b0.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b0.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b0.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b0.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b0.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b0.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b0.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b0.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b0.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b0.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b0.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b0.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b0.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b0.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b0.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b0.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b0.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b0.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b0.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b1.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b1.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b1.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b1.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b1.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b1.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b1.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b1.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b1.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b1.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b1.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b1.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b1.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b1.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b1.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b1.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b1.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b1.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b1.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b1.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b1.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b1.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b1.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b1.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b1.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b1.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b1.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b1.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b1.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b1.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b1.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b1.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b1.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b2.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b2.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b2.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b2.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b2.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b2.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b2.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b2.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b2.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b2.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b2.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b2.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b2.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b2.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b2.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b2.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b2.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b2.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b2.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b2.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b2.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b2.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b2.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b2.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b2.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b2.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b2.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b2.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b2.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b2.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b2.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b2.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b2.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b3.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b3.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b3.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b3.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b3.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b3.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b3.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b3.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b3.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b3.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b3.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b3.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b3.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b3.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b3.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b3.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b3.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b3.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b3.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b3.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b3.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b3.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b3.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b3.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b3.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b3.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b3.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b3.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b3.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b3.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b3.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b3.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b3.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b4.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b4.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b4.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b4.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b4.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b4.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b4.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b4.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b4.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b4.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b4.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b4.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b4.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b4.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b4.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b4.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b4.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b4.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b4.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b4.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b4.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b4.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b4.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b4.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b4.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b4.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b4.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b4.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b4.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b4.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b4.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b4.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b4.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b5.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b5.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b5.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b5.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b5.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b5.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b5.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b5.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b5.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b5.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b5.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b5.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b5.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b5.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b5.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b5.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b5.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b5.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b5.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b5.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b5.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b5.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b5.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b5.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b5.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b5.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b5.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b5.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b5.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b5.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b5.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b5.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b5.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b6.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b6.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b6.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b6.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b6.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b6.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b6.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b6.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b6.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b6.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b6.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b6.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b6.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b6.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b6.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b6.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b6.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b6.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b6.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b6.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b6.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b6.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b6.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b6.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b6.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b6.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b6.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b6.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b6.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b6.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b6.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b6.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b6.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2b7.clock_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2b7.clock_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2b7.evict.ff_evict_control_regs_slice.d0_0 value=000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2b7.evict.ff_evict_control_regs_slice.d0_0.d = 21'b000000000000000000001;

// instance=tb_top.cpu.l2b7.evict.ff_fb_rw_fail.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.l2b7.evict.ff_fb_rw_fail.d0_0.d = 6'b000001;

// instance=tb_top.cpu.l2b7.evict.ff_mux_select0_2b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b7.evict.ff_mux_select0_2b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b7.evict.ff_mux_select1_2a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b7.evict.ff_mux_select1_2a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b7.evict.ff_mux_select2_1b.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b7.evict.ff_mux_select2_1b.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b7.evict.ff_mux_select3_1a.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b7.evict.ff_mux_select3_1a.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b7.evict.ff_rdma_control_regs_slice.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2b7.evict.ff_rdma_control_regs_slice.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2b7.fb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.fb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.fb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.fb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.fb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.fb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.fb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.fb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.fbd.ff_fb_rw_fail.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2b7.fbd.ff_fb_rw_fail.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2b7.fbd.ff_fillbf_control_reg_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b7.fbd.ff_fillbf_control_reg_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b7.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2b7.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2b7.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2b7.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2b7.rdma_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdma_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.rdma_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdma_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.rdma_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdma_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.rdma_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdma_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.rdmard.ff_sel_l1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdmard.ff_sel_l1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b7.rdmard.ff_sel_l2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdmard.ff_sel_l2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b7.rdmard.ff_sel_r1_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdmard.ff_sel_r1_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b7.rdmard.ff_sel_r2_slice.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdmard.ff_sel_r2_slice.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2b7.rdmard.ff_select_inputs.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2b7.rdmard.ff_select_inputs.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2b7.wb_array1.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.wb_array1.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.wb_array2.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.wb_array2.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.wb_array3.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.wb_array3.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2b7.wb_array4.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2b7.wb_array4.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d0.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d0.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d0.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d0.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d0.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d0.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d0.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d0.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d0.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d0.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d0.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d0.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d0.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d0.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d1.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d1.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d1.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d1.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d1.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d1.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d1.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d1.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d1.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d1.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d1.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d1.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d2.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d2.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d2.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d2.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d2.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d2.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d2.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d2.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d2.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d2.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d2.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d2.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d3.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d3.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d3.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d3.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d3.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d3.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d3.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d3.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d3.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d3.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d3.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d3.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d4.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d4.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d4.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d4.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d4.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d4.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d4.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d4.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d4.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d4.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d4.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d4.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d5.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d5.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d5.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d5.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d5.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d5.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d5.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d5.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d5.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d5.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d5.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d5.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d6.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d6.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d6.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d6.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d6.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d6.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d6.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d6.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d6.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d6.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d6.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d6.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c4.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_00.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_20.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_21.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.l2d_clk_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2d7.l2d_clk_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2d7.l2d_clk_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d7.l2d_clk_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2d7.l2d_clk_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d7.l2d_clk_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2d7.l2d_clk_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2d7.l2d_clk_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2d7.l2d_clk_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2d7.l2d_clk_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2d7.perif_io.ff_fill_clk_en_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.perif_io.ff_fill_clk_en_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2d7.perif_io.ff_pwrsav_ov_stg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2d7.perif_io.ff_pwrsav_ov_stg.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t0.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t0.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t0.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t0.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t0.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t0.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t0.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t0.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t0.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t0.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t0.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t0.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t0.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t0.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t0.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t0.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t0.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t0.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t0.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t0.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t0.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t0.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t0.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t0.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t0.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t0.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t0.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t0.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t0.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t0.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t0.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t0.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t0.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t0.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t0.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t0.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t0.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t0.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t0.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t0.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t0.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t0.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t0.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t0.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t0.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t0.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t0.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t0.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t0.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t0.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t0.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t0.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t0.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t0.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t0.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t0.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t0.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t0.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t0.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t0.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t0.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t0.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t0.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t0.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t0.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t0.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t0.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t0.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t0.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t0.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t0.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t0.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t0.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t0.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t0.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t0.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t0.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t1.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t1.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t1.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t1.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t1.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t1.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t1.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t1.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t1.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t1.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t1.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t1.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t1.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t1.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t1.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t1.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t1.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t1.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t1.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t1.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t1.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t1.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t1.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t1.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t1.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t1.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t1.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t1.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t1.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t1.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t1.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t1.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t1.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t1.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t1.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t1.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t1.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t1.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t1.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t1.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t1.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t1.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t1.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t1.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t1.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t1.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t1.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t1.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t1.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t1.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t1.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t1.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t1.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t1.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t1.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t1.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t1.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t1.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t1.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t1.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t1.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t1.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t1.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t1.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t1.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t1.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t1.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t1.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t1.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t1.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t1.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t1.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t1.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t1.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t1.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t1.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t1.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t1.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t2.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t2.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t2.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t2.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t2.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t2.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t2.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t2.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t2.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t2.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t2.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t2.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t2.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t2.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t2.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t2.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t2.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t2.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t2.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t2.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t2.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t2.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t2.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t2.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t2.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t2.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t2.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t2.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t2.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t2.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t2.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t2.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t2.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t2.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t2.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t2.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t2.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t2.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t2.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t2.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t2.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t2.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t2.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t2.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t2.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t2.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t2.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t2.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t2.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t2.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t2.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t2.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t2.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t2.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t2.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t2.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t2.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t2.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t2.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t2.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t2.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t2.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t2.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t2.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t2.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t2.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t2.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t2.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t2.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t2.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t2.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t2.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t2.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t2.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t2.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t2.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t2.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t2.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t3.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t3.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t3.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t3.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t3.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t3.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t3.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t3.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t3.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t3.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t3.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t3.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t3.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t3.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t3.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t3.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t3.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t3.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t3.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t3.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t3.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t3.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t3.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t3.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t3.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t3.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t3.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t3.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t3.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t3.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t3.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t3.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t3.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t3.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t3.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t3.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t3.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t3.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t3.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t3.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t3.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t3.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t3.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t3.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t3.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t3.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t3.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t3.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t3.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t3.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t3.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t3.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t3.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t3.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t3.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t3.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t3.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t3.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t3.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t3.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t3.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t3.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t3.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t3.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t3.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t3.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t3.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t3.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t3.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t3.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t3.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t3.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t3.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t3.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t3.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t3.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t3.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t3.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t4.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t4.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t4.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t4.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t4.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t4.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t4.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t4.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t4.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t4.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t4.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t4.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t4.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t4.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t4.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t4.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t4.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t4.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t4.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t4.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t4.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t4.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t4.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t4.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t4.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t4.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t4.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t4.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t4.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t4.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t4.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t4.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t4.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t4.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t4.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t4.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t4.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t4.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t4.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t4.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t4.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t4.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t4.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t4.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t4.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t4.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t4.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t4.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t4.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t4.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t4.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t4.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t4.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t4.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t4.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t4.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t4.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t4.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t4.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t4.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t4.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t4.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t4.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t4.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t4.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t4.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t4.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t4.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t4.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t4.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t4.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t4.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t4.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t4.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t4.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t4.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t4.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t4.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t5.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t5.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t5.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t5.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t5.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t5.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t5.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t5.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t5.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t5.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t5.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t5.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t5.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t5.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t5.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t5.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t5.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t5.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t5.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t5.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t5.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t5.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t5.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t5.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t5.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t5.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t5.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t5.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t5.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t5.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t5.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t5.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t5.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t5.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t5.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t5.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t5.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t5.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t5.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t5.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t5.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t5.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t5.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t5.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t5.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t5.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t5.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t5.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t5.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t5.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t5.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t5.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t5.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t5.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t5.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t5.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t5.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t5.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t5.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t5.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t5.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t5.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t5.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t5.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t5.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t5.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t5.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t5.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t5.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t5.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t5.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t5.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t5.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t5.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t5.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t5.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t5.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t5.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t6.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t6.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t6.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t6.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t6.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t6.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t6.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t6.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t6.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t6.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t6.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t6.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t6.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t6.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t6.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t6.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t6.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t6.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t6.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t6.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t6.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t6.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t6.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t6.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t6.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t6.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t6.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t6.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t6.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t6.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t6.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t6.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t6.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t6.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t6.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t6.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t6.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t6.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t6.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t6.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t6.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t6.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t6.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t6.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t6.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t6.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t6.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t6.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t6.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t6.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t6.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t6.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t6.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t6.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t6.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t6.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t6.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t6.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t6.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t6.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t6.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t6.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t6.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t6.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t6.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t6.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t6.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t6.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t6.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t6.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t6.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t6.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t6.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t6.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t6.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t6.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t6.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t6.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t7.arb.ff_arb_decdp_cas1_inst_c3.d0_0 value=0001000 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d = 7'b0001000;

// instance=tb_top.cpu.l2t7.arb.ff_data_ecc_active_c4_dup.d0_0 value=01 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.arb.ff_data_ecc_active_c4_dup.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t7.arb.ff_decdp_camld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_decdp_camld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_decdp_ld_inst_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_decdp_ld_inst_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_dword_mask_c8.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_dword_mask_c8.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t7.arb.ff_ic_hitqual_cam_en_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_ic_hitqual_cam_en_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t7.arb.ff_parerr_gate_c1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_parerr_gate_c1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t7.arb.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_waysel_gate_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_waysel_gate_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_word_lower_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_word_lower_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.ff_word_upper_cmp_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.ff_word_upper_cmp_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arb.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.arb.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.arbadr.ff_mux3_bufsel_px2.d0_0 value=00001100 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbadr.ff_mux3_bufsel_px2.d0_0.d = 8'b00001100;

// instance=tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_1.d0_0 value=111100000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_1.d0_0.d = 12'b111100000000;

// instance=tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_2.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_2.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_3.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_3.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t7.arbadr.ff_ncu_signals.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbadr.ff_ncu_signals.d0_0.d = 5'b01111;

// instance=tb_top.cpu.l2t7.arbdat.ff_col_offset_sel_c2.d0_0 value=0001000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbdat.ff_col_offset_sel_c2.d0_0.d = 10'b0001000001;

// instance=tb_top.cpu.l2t7.arbdat.ff_mbdata_mbist_reg.d0_0 value=10000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbdat.ff_mbdata_mbist_reg.d0_0.d = 38'b10000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t7.arbdec.ff_inst_size_c8.d0_0 value=000000000100000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbdec.ff_inst_size_c8.d0_0.d = 18'b000000000100000000;

// instance=tb_top.cpu.l2t7.arbdec.ff_mbdata_mbist_reg.d0_0 value=1100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.arbdec.ff_mbdata_mbist_reg.d0_0.d = 28'b1100000000000000000000000000;

// instance=tb_top.cpu.l2t7.csreg.ff_mux1_sel_c7.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t7.csreg.ff_mux1_sel_c7.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t7.dc_out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.dc_out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.dc_out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.dc_out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.dc_out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.dc_out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.dc_out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.dc_out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.dc_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.dc_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.dc_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.decc.ff_fame_mbist_flops_0.d0_0 value=00000000000000000000000010000 out=q in=d model=dff 
force tb_top.cpu.l2t7.decc.ff_fame_mbist_flops_0.d0_0.d = 29'b00000000000000000000000010000;

// instance=tb_top.cpu.l2t7.deccck.ff_deccck_muxsel_diag_out_c7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.dirrep.ff_dir_vld_dcd_c4_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dirrep.ff_inval_mask_dcd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t7.dirrep.ff_inval_mask_dcd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t7.dirrep.ff_inval_mask_icd_c4.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t7.dirrep.ff_inval_mask_icd_c4.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t7.dirvec.ff_ncu_signals.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.l2t7.dirvec.ff_ncu_signals.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.l2t7.dirvec.ff_staged_part_bank.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t7.dirvec.ff_staged_part_bank.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t7.dirvec.ff_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.dirvec.ff_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.dmologic.ff_dmo_data_1.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.dmologic.ff_dmo_data_1.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t7.evctag.ff_shifted_index.d0_0 value=0000000000000000000000111001100000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.evctag.ff_shifted_index.d0_0.d = 40'b0000000000000000000000111001100000000000;

// instance=tb_top.cpu.l2t7.fbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.fbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.fbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.filbuf.ff_fb_hit_off_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.ff_fb_hit_off_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.filbuf.ff_fill_entry_num_c2.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.ff_fill_entry_num_c2.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.filbuf.ff_fill_entry_num_c3.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.ff_fill_entry_num_c3.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.filbuf.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.filbuf.ff_l2_rd_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.ff_l2_rd_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.filbuf.ff_l2_rd_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.ff_l2_rd_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.filbuf.ff_l2_rd_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.ff_l2_rd_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.filbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.filbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row0.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row0.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row0.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row0.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row0.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row0.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask0_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask0_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask1_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask1_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask2_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask2_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_0 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_0 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_1 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_1 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_1.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_2 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_2 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_2.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_3 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_3 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_3.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_4 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_4 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_4.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_5 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_5 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_5.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_6 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_6 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_6.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_7 value=1 out=latout in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.inv_mask3_so_7 value=1 out=q in=d model=cl_mc1_scm_msff_lat_4x 
force tb_top.cpu.l2t7.ic_row2.inv_mask3_so_7.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.wr_data0_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row2.wr_data0_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.wr_data1_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row2.wr_data1_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.wr_data2_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row2.wr_data2_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.ic_row2.wr_data3_so_15 value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.l2t7.ic_row2.wr_data3_so_15.d = 1'b1;

// instance=tb_top.cpu.l2t7.iqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t7.iqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t7.iqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t7.iqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t7.iqu.ff_array_wr_ptr_plus1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.iqu.ff_array_wr_ptr_plus1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.iqu.ff_iqu_sel_pcx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.iqu.ff_iqu_sel_pcx.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.iqu.ff_que_cnt_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.iqu.ff_que_cnt_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.iqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.iqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.ique.ff_pcx_l2t_data_c1_2.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.ique.ff_pcx_l2t_data_c1_2.d0_0.d = 66'b100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.l2drpt.ff_all_signals.d0_0 value=100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.l2drpt.ff_all_signals.d0_0.d = 21'b100000000000000000000;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.l2t7.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.mb0.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t7.mb0.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t7.mb2_control.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t7.mb2_control.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t7.mbdata.ff_wdata_1.d0_0 value=0000000000000000000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.mbdata.ff_wdata_1.d0_0.d = 64'b0000000000000000000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.mbist.input_signals_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t7.mbist.input_signals_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.l2t7.mbtag.xx84.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.mbtag.xx84.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.mbtag.xx84.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_fbsel_def_vld_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_fbsel_def_vld_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_idx_c1c2comp_c1_d1.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_l2_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_l2_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mb_hit_off_c1_d1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mb_hit_off_c1_d1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t7.misbuf.ff_mb_write_ptr_c3.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mb_write_ptr_c3.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c4.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c4.d0_0.d = 3'b100;

// instance=tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c5.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c52.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c52.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c6.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c7.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_pick_2_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_pick_2_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad4.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad4.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad5.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad5.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad6.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad6.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad7.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad7.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d = 2'b11;

// instance=tb_top.cpu.l2t7.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.misbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.misbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.oqarray.ff_byte_wen.d0_0 value=11111111111111111111 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqarray.ff_byte_wen.d0_0.d = 20'b11111111111111111111;

// instance=tb_top.cpu.l2t7.oqarray.ff_wdata_72.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqarray.ff_wdata_72.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t7.oqarray.ff_word_wen.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqarray.ff_word_wen.d0_0.d = 4'b1111;

// instance=tb_top.cpu.l2t7.oqu.ff_allow_req_c7.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_allow_req_c7.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t7.oqu.ff_dec_cpu_c52.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_dec_cpu_c52.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.oqu.ff_dec_cpu_c6.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_dec_cpu_c6.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.oqu.ff_dec_cpu_c7.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_dec_cpu_c7.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.oqu.ff_dec_cpuid_c6.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_dec_cpuid_c6.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.l2t7.oqu.ff_diag_def_sel_c8.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_diag_def_sel_c8.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.oqu.ff_mux_vec_sel_c52.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_mux_vec_sel_c52.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t7.oqu.ff_mux_vec_sel_c6.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_mux_vec_sel_c6.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t7.oqu.ff_oq_cnt_minus1_d1.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_oq_cnt_minus1_d1.d0_0.d = 5'b11111;

// instance=tb_top.cpu.l2t7.oqu.ff_oq_cnt_plus1_d1.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.ff_oq_cnt_plus1_d1.d0_0.d = 5'b00001;

// instance=tb_top.cpu.l2t7.oqu.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.oqu.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.oque.ff_data_rtn_d1_1.d0_0 value=100000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.oque.ff_data_rtn_d1_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.oque.ff_mbist_flop.d0_0 value=10000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.oque.ff_mbist_flop.d0_0.d = 41'b10000000000000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.oque.ff_tmp_cpx_data_ca_1.d0_0 value=011111111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t7.oque.ff_tmp_cpx_data_ca_1.d0_0.d = 36'b100000000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.out_col0.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.out_col0.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.out_col1.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.out_col1.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.out_col2.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.out_col2.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.out_col3.ff_lookup_cmp_data.d0_0 value=00010000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.out_col3.ff_lookup_cmp_data.d0_0.d = 20'b00010000000000000000;

// instance=tb_top.cpu.l2t7.rdmat.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.rdmat.ff_rdma_wr_ptr_s2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.rdmat.ff_rdma_wr_ptr_s2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.rdmat.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.rdmat.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.rdmatag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.rdmatag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.rdmatag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.l2t7.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d = 2'b10;

// instance=tb_top.cpu.l2t7.snp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.snp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0 value=00000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d = 32'b00000000000000000000000000000001;

// instance=tb_top.cpu.l2t7.subarray_0.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_0.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.subarray_1.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_1.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.subarray_10.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_10.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.subarray_11.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_11.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.subarray_2.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_2.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.subarray_3.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_3.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.subarray_8.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_8.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.subarray_9.ff_word_wen.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.subarray_9.ff_word_wen.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tag.ff_clk_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tag.ff_clk_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.ff_ff_wr_en_ov.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tag.ff_ff_wr_en_ov.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad0.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad0.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad0.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad0.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad0.bank0.reg_wr_way_b.d0_0 value=01 out=latout in=d model=tisram_msff 
force tb_top.cpu.l2t7.tag.quad0.bank0.reg_wr_way_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.l2t7.tag.quad0.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad0.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad0.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad0.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad1.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad1.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad1.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad1.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad1.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad1.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad1.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad1.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad2.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad2.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad2.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad2.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad2.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad2.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad2.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad2.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad3.bank0.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad3.bank0.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad3.bank0.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad3.bank0.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad3.bank1.reg_way_hit_a0.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad3.bank1.reg_way_hit_a0.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tag.quad3.bank1.reg_way_hit_a1.d0_0 value=0 out=q_l in=d model=msffi 
force tb_top.cpu.l2t7.tag.quad3.bank1.reg_way_hit_a1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagctl.ff_alt_tag_miss_unqual_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagctl.ff_l2_bypass_mode_on.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagctl.ff_l2_bypass_mode_on.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagctl.ff_ld_inst_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagctl.ff_ld_inst_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagctl.ff_prev_wen_c1.d0_0 value=0000000000000011 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagctl.ff_prev_wen_c1.d0_0.d = 16'b0000000000000011;

// instance=tb_top.cpu.l2t7.tagctl.ff_scrub_wr_disable_c9.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagctl.ff_scrub_wr_disable_c9.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagctl.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagctl.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagd.ff_ecc_staging5_8.d0_0 value=100000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagd.ff_ecc_staging5_8.d0_0.d = 27'b100000000000000000000000000;

// instance=tb_top.cpu.l2t7.tagd.ff_piped_vuad0.d0_0 value=0000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagd.ff_piped_vuad0.d0_0.d = 28'b0000000000000000000000000001;

// instance=tb_top.cpu.l2t7.tagdp.ff_dir_quad_way_c3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_dir_quad_way_c3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_quad_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_quad_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_state_quad0.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_state_quad0.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_state_quad1.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_state_quad1.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_state_quad2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_state_quad2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_state_quad3.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_state_quad3.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_way_c3.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_way_c3.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t7.tagdp.ff_lru_way_c3_1.d0_0 value=0000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_lru_way_c3_1.d0_0.d = 16'b0000000000000001;

// instance=tb_top.cpu.l2t7.tagdp.ff_tag_quad0_muxsel_c2.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.tagdp.ff_tag_quad1_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t7.tagdp.ff_tag_quad2_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t7.tagdp.ff_tag_quad3_muxsel_c2.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d = 4'b1000;

// instance=tb_top.cpu.l2t7.tagdp.ff_use_dec_sel_c3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.ff_use_dec_sel_c3.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.tagdp.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.tagdp.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.usaloc.ff_used_alloc_c3.d0_0 value=011111111111111111111111111111111 out=q_l in=d model=msffi_dp 
force tb_top.cpu.l2t7.usaloc.ff_used_alloc_c3.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.usaloc.ff_used_and_alloc_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.usaloc.ff_used_and_alloc_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.vlddir.ff_valid_dirty_rd_c2.d0_0 value=100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.l2t7.vlddir.ff_valid_dirty_rd_c2.d0_0.d = 33'b100000000000000000000000000000000;

// instance=tb_top.cpu.l2t7.vuad.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.vuad.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.vuad.ff_vuaddp_vuad_sel_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.vuadpm.ff_mbist_write_data.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.vuadpm.ff_mbist_write_data.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.l2t7.wbtag.xx62.d0_0 value=1 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.wbtag.xx62.d0_0 value=1 out=q in=d model=scm_msff_lat 
force tb_top.cpu.l2t7.wbtag.xx62.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.wbuf.ff_arb_wbuf_hit_off_c2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.wbuf.ff_l2_bypass_mode_on_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.wbuf.ff_quad0_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_quad0_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.wbuf.ff_quad1_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_quad1_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.wbuf.ff_quad2_state.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_quad2_state.d0_0.d = 4'b0001;

// instance=tb_top.cpu.l2t7.wbuf.ff_quad_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_quad_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t7.wbuf.ff_state.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_state.d0_0.d = 3'b001;

// instance=tb_top.cpu.l2t7.wbuf.ff_wbtag_write_wl_c5.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.ff_wbtag_write_wl_c5.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.l2t7.wbuf.reset_flop.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbuf.reset_flop.d0_0.d = 1'b1;

// instance=tb_top.cpu.l2t7.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.l2t7.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d = 3'b010;

// instance=tb_top.cpu.mcu0.clkgen_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu0.clkgen_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu0.clkgen_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu0.clkgen_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu0.clkgen_dr.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu0.clkgen_dr.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu0.clkgen_dr.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu0.clkgen_dr.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu0.clkgen_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu0.clkgen_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu0.drif.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu0.drif.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu0.drif.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu0.drif.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu0.drif.ff_dal_reg.d0_0 value=01101 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.ff_dal_reg.d0_0.d = 5'b01101;

// instance=tb_top.cpu.mcu0.drif.ff_err_fifo_empty_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.ff_err_fifo_empty_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu0.drif.ff_mem_type.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.ff_mem_type.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu0.drif.ff_ral_reg.d0_0 value=01100 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.ff_ral_reg.d0_0.d = 5'b01100;

// instance=tb_top.cpu.mcu0.drif.ff_sync_frame_req_l.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.ff_sync_frame_req_l.d0_0.d = 3'b111;

// instance=tb_top.cpu.mcu0.drif.ff_time_cntr.d0_0 value=0010010010011011 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.ff_time_cntr.d0_0.d = 16'b0010010010011011;

// instance=tb_top.cpu.mcu0.drif.reqq.woq.ff_io_wdata_sel.d0_0 value=0101 out=q in=d model=dff 
force tb_top.cpu.mcu0.drif.reqq.woq.ff_io_wdata_sel.d0_0.d = 4'b0101;

// instance=tb_top.cpu.mcu0.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.ff_chnl_latency_cntr.d0_0 value=10011011 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_chnl_latency_cntr.d0_0.d = 8'b10011011;

// instance=tb_top.cpu.mcu0.fbdic.ff_config_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_config_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu0.fbdic.ff_crc_sel0.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_crc_sel0.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu0.fbdic.ff_crc_sel1.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_crc_sel1.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu0.fbdic.ff_elect_idle_detect.d0_0 value=1111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_elect_idle_detect.d0_0.d = 28'b1111111111111111111111111111;

// instance=tb_top.cpu.mcu0.fbdic.ff_l0s_stall.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_l0s_stall.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu0.fbdic.ff_polling_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_polling_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu0.fbdic.ff_tclktrain_min_cnt.d0_0 value=0000000011111111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_tclktrain_min_cnt.d0_0.d = 16'b0000000011111111;

// instance=tb_top.cpu.mcu0.fbdic.ff_tclktrain_timeout_cnt.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_tclktrain_timeout_cnt.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.mcu0.fbdic.ff_tdisable_cnt.d0_0 value=1100000000 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_tdisable_cnt.d0_0.d = 10'b1100000000;

// instance=tb_top.cpu.mcu0.fbdic.ff_testing_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_testing_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu0.fbdic.ff_ts_match0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_ts_match0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.ff_ts_match0_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_ts_match0_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu0.fbdic.ff_ts_match1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_ts_match1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.ff_ts_match1_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu0.fbdic.ff_ts_match1_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu0.fbdic.spare20_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu0.fbdic.spare20_flop.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll0.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll0.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll0.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll0.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll1.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll1.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll1.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll1.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll2.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll2.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll2.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll2.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll3.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll3.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll3.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll3.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll4.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll4.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll4.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll4.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll5.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll5.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fbdic.sync_stspll5.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu0.fbdic.sync_stspll5.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu0.fdoklu.ff_idle_lfsr.d0_0 value=000000000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.fdoklu.ff_idle_lfsr.d0_0.d = 12'b000000000001;

// instance=tb_top.cpu.mcu0.fdoklu.ff_link_cnt_eq_0_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu0.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu0.fdout.spare0_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu0.fdout.spare0_flop.d = 1'b1;

// instance=tb_top.cpu.mcu0.l2if0.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if0.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu0.l2if0.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if0.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu0.l2if0.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if0.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu0.l2if0.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if0.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu0.l2if0.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if0.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu0.l2if0.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if0.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu0.l2if0.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if0.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu0.l2if1.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu0.l2if1.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu0.l2if1.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu0.l2if1.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu0.l2if1.ff_addr.d0_0 value=00000000000000000000000000000000010 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.ff_addr.d0_0.d = 35'b00000000000000000000000000000000010;

// instance=tb_top.cpu.mcu0.l2if1.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu0.l2if1.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu0.l2if1.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2if1.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu0.l2rdmx.u_l2ecc_mbist_wdata.d0_0 value=0000000000000000000000000000000000000000000000000000001010101011 out=q in=d model=dff 
force tb_top.cpu.mcu0.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d = 64'b0000000000000000000000000000000000000000000000000000001010101011;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw0.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.lndskw1.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu0.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu0.mbist.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu0.mbist.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu0.mbist.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu0.mbist.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu0.mbist.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu0.mbist.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu0.mbist.data_pipe_reg4.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu0.mbist.data_pipe_reg4.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu0.mbist.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu0.mbist.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu0.rdata.ff_ddr_cmp_sync_en_d12.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu0.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu0.rdata.ff_ddr_cmp_sync_en_d23.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu0.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu0.rdata.ff_io_sync_pulses.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu0.rdata.ff_io_sync_pulses.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu0.rdata.ff_mbist_data.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu0.rdata.ff_mbist_data.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.mcu0.rdata.ff_mcu_sync_pulse_delays.d0_0 value=0100 out=q in=d model=dff 
force tb_top.cpu.mcu0.rdata.ff_mcu_sync_pulse_delays.d0_0.d = 4'b0100;

// instance=tb_top.cpu.mcu0.rdata.ff_mcu_sync_pulses.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu0.rdata.ff_mcu_sync_pulses.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu0.rdata.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu0.rdata.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu0.ucb.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu0.ucb.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu0.wrdp.u_io_ecc_15_0.d0_0 value=11110000000000010000000000000000 out=q in=d model=dff 
force tb_top.cpu.mcu0.wrdp.u_io_ecc_15_0.d0_0.d = 32'b11110000000000010000000000000000;

// instance=tb_top.cpu.mcu1.clkgen_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu1.clkgen_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu1.clkgen_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu1.clkgen_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu1.clkgen_dr.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu1.clkgen_dr.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu1.clkgen_dr.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu1.clkgen_dr.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu1.clkgen_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu1.clkgen_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu1.drif.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu1.drif.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu1.drif.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu1.drif.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu1.drif.ff_dal_reg.d0_0 value=01101 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.ff_dal_reg.d0_0.d = 5'b01101;

// instance=tb_top.cpu.mcu1.drif.ff_err_fifo_empty_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.ff_err_fifo_empty_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu1.drif.ff_mem_type.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.ff_mem_type.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu1.drif.ff_ral_reg.d0_0 value=01100 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.ff_ral_reg.d0_0.d = 5'b01100;

// instance=tb_top.cpu.mcu1.drif.ff_sync_frame_req_l.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.ff_sync_frame_req_l.d0_0.d = 3'b111;

// instance=tb_top.cpu.mcu1.drif.ff_time_cntr.d0_0 value=0010010010011001 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.ff_time_cntr.d0_0.d = 16'b0010010010011001;

// instance=tb_top.cpu.mcu1.drif.reqq.woq.ff_io_wdata_sel.d0_0 value=0101 out=q in=d model=dff 
force tb_top.cpu.mcu1.drif.reqq.woq.ff_io_wdata_sel.d0_0.d = 4'b0101;

// instance=tb_top.cpu.mcu1.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.ff_chnl_latency_cntr.d0_0 value=10011001 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_chnl_latency_cntr.d0_0.d = 8'b10011001;

// instance=tb_top.cpu.mcu1.fbdic.ff_config_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_config_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu1.fbdic.ff_crc_sel0.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_crc_sel0.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu1.fbdic.ff_crc_sel1.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_crc_sel1.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu1.fbdic.ff_elect_idle_detect.d0_0 value=1111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_elect_idle_detect.d0_0.d = 28'b1111111111111111111111111111;

// instance=tb_top.cpu.mcu1.fbdic.ff_l0s_stall.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_l0s_stall.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu1.fbdic.ff_polling_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_polling_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu1.fbdic.ff_tclktrain_min_cnt.d0_0 value=0000000011111111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_tclktrain_min_cnt.d0_0.d = 16'b0000000011111111;

// instance=tb_top.cpu.mcu1.fbdic.ff_tclktrain_timeout_cnt.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_tclktrain_timeout_cnt.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.mcu1.fbdic.ff_tdisable_cnt.d0_0 value=1100000000 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_tdisable_cnt.d0_0.d = 10'b1100000000;

// instance=tb_top.cpu.mcu1.fbdic.ff_testing_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_testing_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu1.fbdic.ff_ts_match0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_ts_match0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.ff_ts_match0_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_ts_match0_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu1.fbdic.ff_ts_match1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_ts_match1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.ff_ts_match1_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu1.fbdic.ff_ts_match1_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu1.fbdic.spare20_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu1.fbdic.spare20_flop.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll0.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll0.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll0.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll0.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll1.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll1.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll1.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll1.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll2.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll2.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll2.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll2.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll3.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll3.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll3.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll3.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll4.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll4.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll4.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll4.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll5.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll5.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fbdic.sync_stspll5.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu1.fbdic.sync_stspll5.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu1.fdoklu.ff_idle_lfsr.d0_0 value=000000000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.fdoklu.ff_idle_lfsr.d0_0.d = 12'b000000000001;

// instance=tb_top.cpu.mcu1.fdoklu.ff_link_cnt_eq_0_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu1.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu1.fdout.spare0_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu1.fdout.spare0_flop.d = 1'b1;

// instance=tb_top.cpu.mcu1.l2if0.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if0.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu1.l2if0.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if0.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu1.l2if0.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if0.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu1.l2if0.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if0.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu1.l2if0.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if0.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu1.l2if0.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if0.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu1.l2if0.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if0.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu1.l2if1.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu1.l2if1.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu1.l2if1.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu1.l2if1.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu1.l2if1.ff_addr.d0_0 value=00000000000000000000000000000000010 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.ff_addr.d0_0.d = 35'b00000000000000000000000000000000010;

// instance=tb_top.cpu.mcu1.l2if1.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu1.l2if1.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu1.l2if1.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2if1.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu1.l2rdmx.u_l2ecc_mbist_wdata.d0_0 value=0000000000000000000000000000000000000000000000000000001010101011 out=q in=d model=dff 
force tb_top.cpu.mcu1.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d = 64'b0000000000000000000000000000000000000000000000000000001010101011;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw0.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.lndskw1.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu1.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu1.mbist.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu1.mbist.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu1.mbist.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu1.mbist.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu1.mbist.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu1.mbist.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu1.mbist.data_pipe_reg4.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu1.mbist.data_pipe_reg4.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu1.mbist.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu1.mbist.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu1.rdata.ff_ddr_cmp_sync_en_d12.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu1.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu1.rdata.ff_ddr_cmp_sync_en_d23.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu1.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu1.rdata.ff_io_sync_pulses.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu1.rdata.ff_io_sync_pulses.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu1.rdata.ff_mbist_data.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu1.rdata.ff_mbist_data.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.mcu1.rdata.ff_mcu_sync_pulse_delays.d0_0 value=0100 out=q in=d model=dff 
force tb_top.cpu.mcu1.rdata.ff_mcu_sync_pulse_delays.d0_0.d = 4'b0100;

// instance=tb_top.cpu.mcu1.rdata.ff_mcu_sync_pulses.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu1.rdata.ff_mcu_sync_pulses.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu1.rdata.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu1.rdata.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu1.ucb.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu1.ucb.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu1.wrdp.u_io_ecc_15_0.d0_0 value=11110000000000010000000000000000 out=q in=d model=dff 
force tb_top.cpu.mcu1.wrdp.u_io_ecc_15_0.d0_0.d = 32'b11110000000000010000000000000000;

// instance=tb_top.cpu.mcu2.clkgen_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu2.clkgen_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu2.clkgen_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu2.clkgen_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu2.clkgen_dr.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu2.clkgen_dr.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu2.clkgen_dr.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu2.clkgen_dr.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu2.clkgen_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu2.clkgen_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu2.drif.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu2.drif.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu2.drif.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu2.drif.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu2.drif.ff_dal_reg.d0_0 value=01101 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.ff_dal_reg.d0_0.d = 5'b01101;

// instance=tb_top.cpu.mcu2.drif.ff_err_fifo_empty_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.ff_err_fifo_empty_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu2.drif.ff_mem_type.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.ff_mem_type.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu2.drif.ff_ral_reg.d0_0 value=01100 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.ff_ral_reg.d0_0.d = 5'b01100;

// instance=tb_top.cpu.mcu2.drif.ff_sync_frame_req_l.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.ff_sync_frame_req_l.d0_0.d = 3'b111;

// instance=tb_top.cpu.mcu2.drif.ff_time_cntr.d0_0 value=0010010010010111 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.ff_time_cntr.d0_0.d = 16'b0010010010010111;

// instance=tb_top.cpu.mcu2.drif.reqq.woq.ff_io_wdata_sel.d0_0 value=0101 out=q in=d model=dff 
force tb_top.cpu.mcu2.drif.reqq.woq.ff_io_wdata_sel.d0_0.d = 4'b0101;

// instance=tb_top.cpu.mcu2.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.ff_chnl_latency_cntr.d0_0 value=10010111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_chnl_latency_cntr.d0_0.d = 8'b10010111;

// instance=tb_top.cpu.mcu2.fbdic.ff_config_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_config_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu2.fbdic.ff_crc_sel0.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_crc_sel0.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu2.fbdic.ff_crc_sel1.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_crc_sel1.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu2.fbdic.ff_elect_idle_detect.d0_0 value=1111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_elect_idle_detect.d0_0.d = 28'b1111111111111111111111111111;

// instance=tb_top.cpu.mcu2.fbdic.ff_l0s_stall.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_l0s_stall.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu2.fbdic.ff_polling_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_polling_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu2.fbdic.ff_tclktrain_min_cnt.d0_0 value=0000000011111111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_tclktrain_min_cnt.d0_0.d = 16'b0000000011111111;

// instance=tb_top.cpu.mcu2.fbdic.ff_tclktrain_timeout_cnt.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_tclktrain_timeout_cnt.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.mcu2.fbdic.ff_tdisable_cnt.d0_0 value=1100000000 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_tdisable_cnt.d0_0.d = 10'b1100000000;

// instance=tb_top.cpu.mcu2.fbdic.ff_testing_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_testing_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu2.fbdic.ff_ts_match0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_ts_match0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.ff_ts_match0_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_ts_match0_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu2.fbdic.ff_ts_match1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_ts_match1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.ff_ts_match1_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu2.fbdic.ff_ts_match1_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu2.fbdic.spare20_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu2.fbdic.spare20_flop.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll0.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll0.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll0.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll0.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll1.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll1.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll1.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll1.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll2.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll2.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll2.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll2.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll3.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll3.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll3.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll3.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll4.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll4.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll4.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll4.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll5.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll5.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fbdic.sync_stspll5.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu2.fbdic.sync_stspll5.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu2.fdoklu.ff_idle_lfsr.d0_0 value=000000000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.fdoklu.ff_idle_lfsr.d0_0.d = 12'b000000000001;

// instance=tb_top.cpu.mcu2.fdoklu.ff_link_cnt_eq_0_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu2.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu2.fdout.spare0_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu2.fdout.spare0_flop.d = 1'b1;

// instance=tb_top.cpu.mcu2.l2if0.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if0.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu2.l2if0.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if0.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu2.l2if0.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if0.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu2.l2if0.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if0.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu2.l2if0.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if0.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu2.l2if0.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if0.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu2.l2if0.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if0.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu2.l2if1.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu2.l2if1.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu2.l2if1.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu2.l2if1.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu2.l2if1.ff_addr.d0_0 value=00000000000000000000000000000000010 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.ff_addr.d0_0.d = 35'b00000000000000000000000000000000010;

// instance=tb_top.cpu.mcu2.l2if1.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu2.l2if1.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu2.l2if1.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2if1.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu2.l2rdmx.u_l2ecc_mbist_wdata.d0_0 value=0000000000000000000000000000000000000000000000000000001010101011 out=q in=d model=dff 
force tb_top.cpu.mcu2.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d = 64'b0000000000000000000000000000000000000000000000000000001010101011;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw0.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.lndskw1.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu2.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu2.mbist.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu2.mbist.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu2.mbist.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu2.mbist.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu2.mbist.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu2.mbist.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu2.mbist.data_pipe_reg4.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu2.mbist.data_pipe_reg4.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu2.mbist.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu2.mbist.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu2.rdata.ff_ddr_cmp_sync_en_d12.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu2.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu2.rdata.ff_ddr_cmp_sync_en_d23.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu2.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu2.rdata.ff_io_sync_pulses.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu2.rdata.ff_io_sync_pulses.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu2.rdata.ff_mbist_data.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu2.rdata.ff_mbist_data.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.mcu2.rdata.ff_mcu_sync_pulse_delays.d0_0 value=0100 out=q in=d model=dff 
force tb_top.cpu.mcu2.rdata.ff_mcu_sync_pulse_delays.d0_0.d = 4'b0100;

// instance=tb_top.cpu.mcu2.rdata.ff_mcu_sync_pulses.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu2.rdata.ff_mcu_sync_pulses.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu2.rdata.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu2.rdata.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu2.ucb.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu2.ucb.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu2.wrdp.u_io_ecc_15_0.d0_0 value=11110000000000010000000000000000 out=q in=d model=dff 
force tb_top.cpu.mcu2.wrdp.u_io_ecc_15_0.d0_0.d = 32'b11110000000000010000000000000000;

// instance=tb_top.cpu.mcu3.clkgen_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu3.clkgen_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu3.clkgen_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu3.clkgen_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu3.clkgen_dr.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mcu3.clkgen_dr.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mcu3.clkgen_dr.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu3.clkgen_dr.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu3.clkgen_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mcu3.clkgen_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mcu3.drif.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu3.drif.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu3.drif.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu3.drif.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu3.drif.ff_dal_reg.d0_0 value=01101 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.ff_dal_reg.d0_0.d = 5'b01101;

// instance=tb_top.cpu.mcu3.drif.ff_err_fifo_empty_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.ff_err_fifo_empty_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu3.drif.ff_mem_type.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.ff_mem_type.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu3.drif.ff_ral_reg.d0_0 value=01100 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.ff_ral_reg.d0_0.d = 5'b01100;

// instance=tb_top.cpu.mcu3.drif.ff_sync_frame_req_l.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.ff_sync_frame_req_l.d0_0.d = 3'b111;

// instance=tb_top.cpu.mcu3.drif.ff_time_cntr.d0_0 value=0010010010010101 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.ff_time_cntr.d0_0.d = 16'b0010010010010101;

// instance=tb_top.cpu.mcu3.drif.reqq.woq.ff_io_wdata_sel.d0_0 value=0101 out=q in=d model=dff 
force tb_top.cpu.mcu3.drif.reqq.woq.ff_io_wdata_sel.d0_0.d = 4'b0101;

// instance=tb_top.cpu.mcu3.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.ff_chnl_latency_cntr.d0_0 value=10010101 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_chnl_latency_cntr.d0_0.d = 8'b10010101;

// instance=tb_top.cpu.mcu3.fbdic.ff_config_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_config_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu3.fbdic.ff_crc_sel0.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_crc_sel0.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu3.fbdic.ff_crc_sel1.d0_0 value=10100 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_crc_sel1.d0_0.d = 5'b10100;

// instance=tb_top.cpu.mcu3.fbdic.ff_elect_idle_detect.d0_0 value=1111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_elect_idle_detect.d0_0.d = 28'b1111111111111111111111111111;

// instance=tb_top.cpu.mcu3.fbdic.ff_l0s_stall.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_l0s_stall.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu3.fbdic.ff_polling_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_polling_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu3.fbdic.ff_tclktrain_min_cnt.d0_0 value=0000000011111111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_tclktrain_min_cnt.d0_0.d = 16'b0000000011111111;

// instance=tb_top.cpu.mcu3.fbdic.ff_tclktrain_timeout_cnt.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_tclktrain_timeout_cnt.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.mcu3.fbdic.ff_tdisable_cnt.d0_0 value=1100000000 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_tdisable_cnt.d0_0.d = 10'b1100000000;

// instance=tb_top.cpu.mcu3.fbdic.ff_testing_timeout_cnt.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_testing_timeout_cnt.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.mcu3.fbdic.ff_ts_match0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_ts_match0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.ff_ts_match0_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_ts_match0_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu3.fbdic.ff_ts_match1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_ts_match1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.ff_ts_match1_cnt.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.mcu3.fbdic.ff_ts_match1_cnt.d0_0.d = 4'b1111;

// instance=tb_top.cpu.mcu3.fbdic.spare20_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu3.fbdic.spare20_flop.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll0.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll0.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll0.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll0.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll1.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll1.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll1.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll1.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll2.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll2.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll2.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll2.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll3.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll3.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll3.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll3.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll4.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll4.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll4.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll4.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll5.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll5.xx0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fbdic.sync_stspll5.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mcu3.fbdic.sync_stspll5.xx1.d = 1'b1;

// instance=tb_top.cpu.mcu3.fdoklu.ff_idle_lfsr.d0_0 value=000000000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.fdoklu.ff_idle_lfsr.d0_0.d = 12'b000000000001;

// instance=tb_top.cpu.mcu3.fdoklu.ff_link_cnt_eq_0_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu3.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu3.fdout.spare0_flop value=1 out=q in=d model=cl_sc1_msff_8x 
force tb_top.cpu.mcu3.fdout.spare0_flop.d = 1'b1;

// instance=tb_top.cpu.mcu3.l2if0.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if0.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu3.l2if0.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if0.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu3.l2if0.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if0.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu3.l2if0.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if0.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu3.l2if0.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if0.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu3.l2if0.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if0.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu3.l2if0.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if0.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu3.l2if1.adrgen.ff_error_mask.d0_0 value=1111000 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.adrgen.ff_error_mask.d0_0.d = 7'b1111000;

// instance=tb_top.cpu.mcu3.l2if1.adrgen.ff_mem_type.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.adrgen.ff_mem_type.d0_0.d = 4'b1000;

// instance=tb_top.cpu.mcu3.l2if1.adrgen.ff_num_dimms.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.adrgen.ff_num_dimms.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.mcu3.l2if1.adrgen.ff_rank_mask.d0_0 value=000000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.adrgen.ff_rank_mask.d0_0.d = 9'b000000001;

// instance=tb_top.cpu.mcu3.l2if1.ff_addr.d0_0 value=00000000000000000000000000000000010 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.ff_addr.d0_0.d = 35'b00000000000000000000000000000000010;

// instance=tb_top.cpu.mcu3.l2if1.ff_addr_mode.d0_0 value=00110010 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.ff_addr_mode.d0_0.d = 8'b00110010;

// instance=tb_top.cpu.mcu3.l2if1.ff_mcu_sync_pulses.d0_0 value=110 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.ff_mcu_sync_pulses.d0_0.d = 3'b110;

// instance=tb_top.cpu.mcu3.l2if1.ff_partial_mode.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2if1.ff_partial_mode.d0_0.d = 3'b100;

// instance=tb_top.cpu.mcu3.l2rdmx.u_l2ecc_mbist_wdata.d0_0 value=0000000000000000000000000000000000000000000000000000001010101011 out=q in=d model=dff 
force tb_top.cpu.mcu3.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d = 64'b0000000000000000000000000000000000000000000000000000001010101011;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw0.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf0.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf1.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf10.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf11.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf12.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf13.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf2.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf3.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf4.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf5.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf6.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf7.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf8.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.lndskw1.algnbf9.ff_rptr_wptr.d0_0 value=000001 out=q in=d model=dff 
force tb_top.cpu.mcu3.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d = 6'b000001;

// instance=tb_top.cpu.mcu3.mbist.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu3.mbist.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu3.mbist.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu3.mbist.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu3.mbist.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu3.mbist.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu3.mbist.data_pipe_reg4.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu3.mbist.data_pipe_reg4.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu3.mbist.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.mcu3.mbist.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.mcu3.rdata.ff_ddr_cmp_sync_en_d12.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu3.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu3.rdata.ff_ddr_cmp_sync_en_d23.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.mcu3.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d = 1'b1;

// instance=tb_top.cpu.mcu3.rdata.ff_io_sync_pulses.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.mcu3.rdata.ff_io_sync_pulses.d0_0.d = 2'b10;

// instance=tb_top.cpu.mcu3.rdata.ff_mbist_data.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.mcu3.rdata.ff_mbist_data.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.mcu3.rdata.ff_mcu_sync_pulse_delays.d0_0 value=0100 out=q in=d model=dff 
force tb_top.cpu.mcu3.rdata.ff_mcu_sync_pulse_delays.d0_0.d = 4'b0100;

// instance=tb_top.cpu.mcu3.rdata.ff_mcu_sync_pulses.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.mcu3.rdata.ff_mcu_sync_pulses.d0_0.d = 2'b11;

// instance=tb_top.cpu.mcu3.rdata.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu3.rdata.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu3.ucb.ff_partial_bank_mode.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.mcu3.ucb.ff_partial_bank_mode.d0_0.d = 5'b01111;

// instance=tb_top.cpu.mcu3.wrdp.u_io_ecc_15_0.d0_0 value=11110000000000010000000000000000 out=q in=d model=dff 
force tb_top.cpu.mcu3.wrdp.u_io_ecc_15_0.d0_0.d = 32'b11110000000000010000000000000000;

// instance=tb_top.cpu.mio.cell_10.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_10.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_103.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_103.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_104.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_104.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_105.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_105.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_106.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_106.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_107.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_107.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_108.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_108.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_110.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_110.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_12.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_12.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_129.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_129.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_13.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_13.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_130.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_130.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_131.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_131.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_132.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_132.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_133.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_133.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_134.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_134.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_135.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_135.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_136.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_136.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_137.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_137.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_138.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_138.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_139.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_139.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_14.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_14.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_140.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_140.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_141.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_141.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_142.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_142.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_143.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_143.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_144.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_144.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_145.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_145.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_146.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_146.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_147.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_147.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_148.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_148.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_149.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_149.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_15.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_15.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_15.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_15.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_150.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_150.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_151.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_151.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_152.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_152.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_153.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_153.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_154.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_154.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_155.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_155.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_156.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_156.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_157.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_157.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_158.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_158.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_159.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_159.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_160.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_160.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_161.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_161.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_162.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_162.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_163.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_163.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_164.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_164.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_165.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_165.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_17.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_17.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_176.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_176.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_177.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_177.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_178.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_178.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_179.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_179.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_18.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_18.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_180.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_180.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_181.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_181.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_182.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_182.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_184.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_184.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_186.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_186.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_187.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_187.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_189.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_189.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_193.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_193.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_2.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_2.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_202.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_202.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_209.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_209.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_210.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_210.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_211.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_211.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_211.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_211.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_23.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_23.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_24.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_24.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_27.ff_in_mux_data.d0_0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mio.cell_27.ff_in_mux_data.d0_0.d = 1'b1;

// instance=tb_top.cpu.mio.cell_3.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_3.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_3.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_3.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_4.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_4.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.cell_5.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_5.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_6.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_6.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_7.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_7.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_7.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_7.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_8.ff_in value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_8.ff_in.d = 1'b1;

// instance=tb_top.cpu.mio.cell_9.ff_oe value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_9.ff_oe.d = 1'b1;

// instance=tb_top.cpu.mio.cell_9.ff_out value=1 out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_9.ff_out.d = 1'b1;

// instance=tb_top.cpu.mio.cell_98.ff_in value=z out=q in=d model=cl_sc1_bs_cell2_4x 
force tb_top.cpu.mio.cell_98.ff_in.d = 1'bz;

// instance=tb_top.cpu.mio.io2xsyncen_reg0.ff_0.d0_0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mio.io2xsyncen_reg0.ff_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mio.io2xsyncen_reg1.ff_0.d0_0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mio.io2xsyncen_reg1.ff_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mio.io2xsyncen_reg2.ff_0.d0_0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mio.io2xsyncen_reg2.ff_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mio.io2xsyncen_reg3.ff_0.d0_0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mio.io2xsyncen_reg3.ff_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.mio.mio_clk_header_iol2clk.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.mio.mio_clk_header_iol2clk.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.mio.muxsel.ff_1.d0_1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.mio.muxsel.ff_1.d0_1.d = 1'b1;

// instance=tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.ncu.clkgen_ncu_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.ncu.clkgen_ncu_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_cpu_buf_rf_cust.dff_din_hi.d0_0 value=111111111100000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_cpu_buf_rf_cust.dff_din_hi.d0_0.d = 72'b111111111100000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_cpu_buf_rf_cust.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_cpu_buf_rf_cust.dff_dout.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_din_hi.d0_0 value=111111111111101100000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_din_hi.d0_0.d = 72'b111111111111101100000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_din_lo.d0_0 value=000000000000000000000000000000000000000000000000000000000000000000000100 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_din_lo.d0_0.d = 72'b000000000000000000000000000000000000000000000000000000000000000000000100;

// instance=tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_dout.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_din_hi.d0_0 value=111111111111101100000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_din_hi.d0_0.d = 72'b111111111111101100000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_din_lo.d0_0 value=000000000000000000000000000000000000000000000000000000000000000000000100 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_din_lo.d0_0.d = 72'b000000000000000000000000000000000000000000000000000000000000000000000100;

// instance=tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_dout.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.io_cmp_sync_en_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.io_cmp_sync_en_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifc_ctl.cpu_mondo_addr_creg_mdata0_dec_d1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifc_ctl.cpu_mondo_addr_creg_mdata0_dec_d1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo2cpu_pkt_ff.d0_0 value=00000001101000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo2cpu_pkt_ff.d0_0.d = 122'b00000001101000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_busy_dout_d2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_busy_dout_d2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_busy_vec_ff.d0_0 value=1111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_busy_vec_ff.d0_0.d = 64'b1111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data0_din_d1_ff.d0_0 value=111111110000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data0_din_d1_ff.d0_0.d = 72'b111111110000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data0_din_d2_ff.d0_0 value=111111110000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data0_din_d2_ff.d0_0.d = 72'b111111110000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data1_din_d1_ff.d0_0 value=111111110000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data1_din_d1_ff.d0_0.d = 72'b111111110000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data1_din_d2_ff.d0_0 value=111111110000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data1_din_d2_ff.d0_0.d = 72'b111111110000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.intbuf_pa_ff.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.intbuf_pa_ff.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.iobuf_pa_ff.d0_0 value=11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.iobuf_pa_ff.d0_0.d = 176'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.mb0_wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.mb0_wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.res_read_data_reg.d0_0 value=111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.res_read_data_reg.d0_0.d = 48'b111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_intbuf_rf_cust.dff_din_hi.d0_0 value=011111111010111110011100000001101000001000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_intbuf_rf_cust.dff_din_hi.d0_0.d = 72'b011111111010111110011100000001101000001000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_intbuf_rf_cust.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_intbuf_rf_cust.dff_dout.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_intman_rf_cust.dff_din_hi.d0_0 value=11110000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_intman_rf_cust.dff_din_hi.d0_0.d = 8'b11110000;

// instance=tb_top.cpu.ncu.ncu_intman_rf_cust.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.ncu.ncu_intman_rf_cust.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_intman_rf_cust.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.ncu.ncu_intman_rf_cust.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_iobuf0_rf_cust.dff_din_hi.d0_0 value=000010100000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_iobuf0_rf_cust.dff_din_hi.d0_0.d = 72'b000010100000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_iobuf0_rf_cust.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_iobuf0_rf_cust.dff_dout.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_din_hi.d0_0 value=1001111010111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_din_hi.d0_0.d = 16'b1001111010111111;

// instance=tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_din_lo.d0_0 value=1100111000000011 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_din_lo.d0_0.d = 16'b1100111000000011;

// instance=tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_dout.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_dout.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_din_hi.d0_0 value=111111110000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_din_hi.d0_0.d = 36'b111111110000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_din_hi.d0_0 value=111111110000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_din_hi.d0_0.d = 36'b111111110000000000000000000000000000;

// instance=tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ccu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ccu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ccu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ccu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dbg1_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dbg1_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dbg1_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dbg1_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmucsr_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmucsr_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmucsr_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmucsr_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.cr_id_rtn1_par_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.cr_id_rtn1_par_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.ncu_dmu_dpar_ff.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.ncu_dmu_dpar_ff.d0_0.d = 2'b11;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.pad_ff.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.pad_ff.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu0_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu0_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu0_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu0_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu1_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu1_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu1_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu1_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu2_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu2_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu2_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu2_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu3_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu3_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu3_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu3_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_c2isd_ctl.cpubuf_pa_ff.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_c2isd_ctl.cpubuf_pa_ff.d0_0.d = 144'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.core_running_status0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.core_running_status0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.fusestat_ff.d0_0 value=1111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.fusestat_ff.d0_0.d = 64'b1111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.l2pm_ff.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.l2pm_ff.d0_0.d = 5'b01111;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.l2pm_preview_ff.d0_0 value=11111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.l2pm_preview_ff.d0_0.d = 5'b11111;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.por_upd_en_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.por_upd_en_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg1.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg1.d0_0.d = 2'b11;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg2.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg2.d0_0.d = 2'b11;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg3.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg3.d0_0.d = 2'b11;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg4.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg4.d0_0.d = 2'b11;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.mb1_wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.mb1_wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.res_read_data_reg.d0_0 value=1111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.res_read_data_reg.d0_0.d = 40'b1111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.niu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.niu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.niu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.niu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.rcu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.rcu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.rcu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.rcu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ssi_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ssi_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ssi_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ssi_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.tcu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.tcu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.tcu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.tcu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ccu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ccu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ccu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ccu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dbg1_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dbg1_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dbg1_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dbg1_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dmucsr_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dmucsr_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dmucsr_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dmucsr_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu0_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu0_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu0_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu0_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu1_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu1_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu1_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu1_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu2_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu2_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu2_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu2_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu3_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu3_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu3_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu3_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ncu_i2csc_ctl.mondo_busy_d1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ncu_i2csc_ctl.mondo_busy_d1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ncu_i2csc_ctl.mondo_busy_vec_ff.d0_0 value=1111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ncu_i2csc_ctl.mondo_busy_vec_ff.d0_0.d = 64'b1111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.niu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.niu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.niu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.niu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.rcu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.rcu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.rcu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.rcu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.ncu_dmu_mondo_id_par_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.ncu_dmu_mondo_id_par_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ssi_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ssi_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ssi_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ssi_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.tcu_ucb_buf.rdy0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.tcu_ucb_buf.rdy0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.tcu_ucb_buf.rdy1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.tcu_ucb_buf.rdy1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.cntr_ff.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.cntr_ff.d0_0.d = 3'b111;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.sck_cnt_ff.d0_0 value=000000001001001001 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.sck_cnt_ff.d0_0.d = 18'b000000001001001001;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.sck_posedge_d3_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.sck_posedge_d3_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_async_ctu_jbi_ssiclk_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_async_ctu_jbi_ssiclk_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_async_jbi_io_ssi_sck.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_async_jbi_io_ssi_sck.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_sck_cyc_cnt.d0_0 value=1001001 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_sck_cyc_cnt.d0_0.d = 7'b1001001;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg3.p_out_ff.d0_0 value=11000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg3.p_out_ff.d0_0.d = 8'b11000000;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg4.p_out_ff.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg4.p_out_ff.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg5.p_out_ff.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg5.p_out_ff.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg6.p_out_ff.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg6.p_out_ff.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg7.p_out_ff.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg7.p_out_ff.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.toreg_ld0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.toreg_ld0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.toreg_ld1_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.toreg_ld1_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d1.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d2.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d2.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d3.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d3.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d4.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d4.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d5.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d5.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d6.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d6.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d7.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d7.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_io_jbi_ext_int_l_pre_sync.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_io_jbi_ext_int_l_pre_sync.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_io_jbi_ext_int_l_sync.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_io_jbi_ext_int_l_sync.d0_0.d = 1'b1;

// instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_timeout_reg.d0_0 value=0001000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_timeout_reg.d0_0.d = 25'b0001000000000000000000000;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.rst.clkgen_rst_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.ccu_rst_change_cmp0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.ccu_rst_change_cmp0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.ccu_rst_change_cmp_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.ccu_rst_change_cmp_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.io_cmp_sync_en2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.io_cmp_sync_en2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.mio_rst_pb_rst_cmp_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.mio_rst_pb_rst_cmp_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.mio_rst_pb_rst_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.mio_rst_pb_rst_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_cmp_ctl_wmr_cmp_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_cmp_ctl_wmr_cmp_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_dmu_peu_por_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_dmu_peu_por_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_dmu_peu_wmr_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_dmu_peu_wmr_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_l2_por_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_l2_por_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_l2_wmr_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_l2_wmr_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_niu_mac_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_niu_mac_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_niu_wmr_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_niu_wmr_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_rst_por_cmp_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_rst_por_cmp_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_rst_por_io_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_rst_por_io_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_rst_pwron_rst_l_io0_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_rst_pwron_rst_l_io0_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_rst_wmr_cmp_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_rst_wmr_cmp_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_rst_wmr_io_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_rst_wmr_io_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.rst_tcu_pwron_rst_l_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.rst_tcu_pwron_rst_l_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_cmp_ctl.tcu_rst_flush_stop_ack_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_cmp_ctl.tcu_rst_flush_stop_ack_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.ccu_count_ff.d0_0 value=0000000000100000 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.ccu_count_ff.d0_0.d = 16'b0000000000100000;

// instance=tb_top.cpu.rst.rst_fsm_ctl.ccu_rst_change_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.ccu_rst_change_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.cluster_arst_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.cluster_arst_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.lock_count_ff.d0_0 value=0000000000010000 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.lock_count_ff.d0_0.d = 16'b0000000000010000;

// instance=tb_top.cpu.rst.rst_fsm_ctl.mio_rst_button_xir_sys_ff.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.rst.rst_fsm_ctl.mio_rst_button_xir_sys_ff.xx0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.mio_rst_button_xir_sys_ff.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.rst.rst_fsm_ctl.mio_rst_button_xir_sys_ff.xx1.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys3_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys3_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys_ff.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys_ff.xx0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys_ff.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys_ff.xx1.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pwron_rst_sys_ff.xx0 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pwron_rst_sys_ff.xx0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pwron_rst_sys_ff.xx1 value=1 out=q in=d model=cl_sc1_msff_4x 
force tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pwron_rst_sys_ff.xx1.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.niu_count_ff.d0_0 value=0000011001000000 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.niu_count_ff.d0_0.d = 16'b0000011001000000;

// instance=tb_top.cpu.rst.rst_fsm_ctl.prop_count_ff.d0_0 value=0000000000010000 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.prop_count_ff.d0_0.d = 16'b0000000000010000;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_ccu_pll_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_ccu_pll_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_ccu_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_ccu_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_cmp_ctl_wmr_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_cmp_ctl_wmr_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_async_por_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_async_por_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_peu_por_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_peu_por_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_peu_wmr_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_peu_wmr_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_l2_por_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_l2_por_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_l2_wmr_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_l2_wmr_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_niu_mac_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_niu_mac_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_niu_wmr_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_niu_wmr_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_rst_por_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_rst_por_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_rst_pwron_rst_sys2_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_rst_pwron_rst_sys2_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.rst_rst_wmr_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.rst_rst_wmr_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_fsm_ctl.state_ff.d0_0 value=000000000000000000000100000000001 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.state_ff.d0_0.d = 33'b000000000000000000000100000000001;

// instance=tb_top.cpu.rst.rst_fsm_ctl.tr_flush_stop_ack_sys_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_fsm_ctl.tr_flush_stop_ack_sys_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_io_ctl.ccu_rst_change_io_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_io_ctl.ccu_rst_change_io_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_io_ctl.rst_rst_por_io_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_io_ctl.rst_rst_por_io_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_io_ctl.rst_rst_pwron_rst_l_io_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_io_ctl.rst_rst_pwron_rst_l_io_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.rst.rst_io_ctl.rst_rst_wmr_io_ff.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.rst.rst_io_ctl.rst_rst_wmr_io_ff.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.clkgen_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.sii.clkgen_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.sii.clkgen_cmp.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.sii.clkgen_cmp.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.sii.clkgen_cmp.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.sii.clkgen_cmp.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.sii.clkgen_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.sii.clkgen_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.sii.clkgen_cmp.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.sii.clkgen_cmp.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.sii.clkgen_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.sii.clkgen_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.sii.clkgen_io.xcluster_header.control_sig_sync.slow_cmp_sync_en_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.sii.clkgen_io.xcluster_header.control_sig_sync.slow_cmp_sync_en_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.sii.ilc0.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc0.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc0.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc0.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc0.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc0.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ilc1.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc1.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc1.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc1.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc1.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc1.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ilc2.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc2.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc2.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc2.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc2.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc2.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ilc3.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc3.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc3.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc3.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc3.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc3.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ilc4.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc4.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc4.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc4.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc4.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc4.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ilc5.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc5.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc5.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc5.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc5.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc5.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ilc6.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc6.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc6.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc6.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc6.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc6.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ilc7.reg_ilc_ild_addr_h.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc7.reg_ilc_ild_addr_h.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc7.reg_ilc_ild_addr_lo.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.sii.ilc7.reg_ilc_ild_addr_lo.d0_0.d = 4'b0001;

// instance=tb_top.cpu.sii.ilc7.reg_ilc_ildq_rd_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ilc7.reg_ilc_ildq_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ild0.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild0.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild1.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild1.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild2.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild2.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild3.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild3.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild4.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild4.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild5.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild5.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild6.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild6.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild7.ff_sii_mb0_ild_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.ild7.ff_sii_mb0_ild_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_r.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_r.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_rr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_rr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_rrr.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_rrr.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ildq0.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq0.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq0.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq0.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq1.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq1.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq1.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq1.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq2.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq2.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq2.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq2.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq3.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq3.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq3.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq3.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq4.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq4.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq4.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq4.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq5.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq5.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq5.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq5.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq6.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq6.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq6.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq6.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq7.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ildq7.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ildq7.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ildq7.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.inc.reg_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.inc.reg_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.inc.reg_mbist1_data_r.d0_0 value=01010101010101010101010101010101010101010101010101010101010101010101 out=q in=d model=dff 
force tb_top.cpu.sii.inc.reg_mbist1_data_r.d0_0.d = 68'b01010101010101010101010101010101010101010101010101010101010101010101;

// instance=tb_top.cpu.sii.inc.reg_mbist1_data_rr.d0_0 value=01010101010101010101010101010101010101010101010101010101010101010101 out=q in=d model=dff 
force tb_top.cpu.sii.inc.reg_mbist1_data_rr.d0_0.d = 68'b01010101010101010101010101010101010101010101010101010101010101010101;

// instance=tb_top.cpu.sii.inc.reg_sii_mb0_ind_fail.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.inc.reg_sii_mb0_ind_fail.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.inc.reg_sii_mb0_wdata.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.inc.reg_sii_mb0_wdata.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.indq.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.indq.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.indq.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.indq.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipcc.reg_arb1.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.sii.ipcc.reg_arb1.d0_0.d = 2'b10;

// instance=tb_top.cpu.sii.ipcc.reg_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ipcc.reg_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipcc.reg_ncu_sii_ba01.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ipcc.reg_ncu_sii_ba01.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipcc.reg_ncu_sii_ba23.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ipcc.reg_ncu_sii_ba23.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipcc.reg_ncu_sii_ba45.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ipcc.reg_ncu_sii_ba45.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipcc.reg_ncu_sii_ba67.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sii.ipcc.reg_ncu_sii_ba67.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipcc_dp.ff_mb0_wdata.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.ipcc_dp.ff_mb0_wdata.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.ipdbdq0_h.dff_din_hi.d0_0 value=0000000011111111000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.sii.ipdbdq0_h.dff_din_hi.d0_0.d = 40'b0000000011111111000000000000000000000000;

// instance=tb_top.cpu.sii.ipdbdq0_h.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq0_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbdq0_h.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq0_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbdq0_l.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq0_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbdq0_l.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq0_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbdq1_h.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq1_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbdq1_h.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq1_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbdq1_l.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq1_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbdq1_l.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdbdq1_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbhq0.dff_din_hi.d0_0 value=000000001001000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.sii.ipdbhq0.dff_din_hi.d0_0.d = 36'b000000001001000000000000000000000000;

// instance=tb_top.cpu.sii.ipdbhq0.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdbhq0.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbhq0.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdbhq0.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbhq1.dff_din_hi.d0_0 value=000000001001000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.sii.ipdbhq1.dff_din_hi.d0_0.d = 36'b000000001001000000000000000000000000;

// instance=tb_top.cpu.sii.ipdbhq1.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdbhq1.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdbhq1.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdbhq1.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq0_h.dff_din_hi.d0_0 value=0000000011111111000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.sii.ipdodq0_h.dff_din_hi.d0_0.d = 40'b0000000011111111000000000000000000000000;

// instance=tb_top.cpu.sii.ipdodq0_h.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq0_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq0_h.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq0_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq0_l.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq0_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq0_l.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq0_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq1_h.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq1_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq1_h.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq1_h.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq1_l.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq1_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdodq1_l.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdodq1_l.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdohq0.dff_din_hi.d0_0 value=000000001001000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.sii.ipdohq0.dff_din_hi.d0_0.d = 36'b000000001001000000000000000000000000;

// instance=tb_top.cpu.sii.ipdohq0.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdohq0.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdohq0.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdohq0.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdohq1.dff_din_hi.d0_0 value=000000001001000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.sii.ipdohq1.dff_din_hi.d0_0.d = 36'b000000001001000000000000000000000000;

// instance=tb_top.cpu.sii.ipdohq1.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.sii.ipdohq1.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.ipdohq1.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.sii.ipdohq1.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sii.mb0.ild0_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild0_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ild1_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild1_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ild2_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild2_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ild3_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild3_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ild4_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild4_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ild5_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild5_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ild6_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild6_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ild7_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ild7_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.ind_fail_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.ind_fail_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.sii.mb0.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb0.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.mb1.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.mb1.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.mb1.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.mb1.data_pipe_reg4.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.data_pipe_reg4.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.mb1.data_pipe_reg5.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.data_pipe_reg5.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.mb1.sel_pipe_reg1.d0_0 value=000100 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.sel_pipe_reg1.d0_0.d = 6'b000100;

// instance=tb_top.cpu.sii.mb1.sel_pipe_reg2.d0_0 value=000100 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.sel_pipe_reg2.d0_0.d = 6'b000100;

// instance=tb_top.cpu.sii.mb1.sel_reg.d0_0 value=000100 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.sel_reg.d0_0.d = 6'b000100;

// instance=tb_top.cpu.sii.mb1.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sii.mb1.wdata_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sii.mb1.wdata_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.clkgen_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.sio.clkgen_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.sio.clkgen_cmp.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.sio.clkgen_cmp.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.sio.clkgen_cmp.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.sio.clkgen_cmp.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.sio.clkgen_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.sio.clkgen_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.sio.clkgen_cmp.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.sio.clkgen_cmp.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.sio.clkgen_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.sio.clkgen_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.sio.clkgen_io.xcluster_header.control_sig_sync.slow_cmp_sync_en_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.sio.clkgen_io.xcluster_header.control_sig_sync.slow_cmp_sync_en_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.sio.mb0.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb0.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb0.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb0.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb0.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb0.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb0.data_pipe_reg4.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb0.data_pipe_reg4.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb0.read_data_pipe_reg.d0_0 value=11111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.mb0.read_data_pipe_reg.d0_0.d = 68'b11111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.mb0.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb0.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb1.data_pipe_reg1.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.data_pipe_reg1.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb1.data_pipe_reg2.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.data_pipe_reg2.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb1.data_pipe_reg3.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.data_pipe_reg3.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.mb1.opd_sel_reg1.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.opd_sel_reg1.d0_0.d = 3'b010;

// instance=tb_top.cpu.sio.mb1.opd_sel_reg2.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.opd_sel_reg2.d0_0.d = 3'b010;

// instance=tb_top.cpu.sio.mb1.opd_sel_reg4.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.opd_sel_reg4.d0_0.d = 3'b010;

// instance=tb_top.cpu.sio.mb1.read_data_pipe_reg.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.read_data_pipe_reg.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.mb1.sel_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.sel_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.sio.mb1.wdata_reg.d0_0 value=01010101 out=q in=d model=dff 
force tb_top.cpu.sio.mb1.wdata_reg.d0_0.d = 8'b01010101;

// instance=tb_top.cpu.sio.olddq00.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq00.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq01.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq01.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq10.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq10.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq11.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq11.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq20.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq20.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq21.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq21.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq30.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq30.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq31.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq31.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq40.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq40.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq41.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq41.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq50.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq50.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq51.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq51.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq60.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq60.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq61.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq61.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq70.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq70.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.olddq71.dff_dout.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.olddq71.dff_dout.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opcc.reg_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sio.opcc.reg_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.sio.opcs0.reg_opdhqx_ue_bit.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sio.opcs0.reg_opdhqx_ue_bit.d0_0.d = 1'b1;

// instance=tb_top.cpu.sio.opcs1.reg_opdhqx_ue_bit.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.sio.opcs1.reg_opdhqx_ue_bit.d0_0.d = 1'b1;

// instance=tb_top.cpu.sio.opdc.dff_bank01_data_opc1_h.d0_0 value=0111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank01_data_opc1_h.d0_0.d = 34'b0111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_bank01_data_opc1_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank01_data_opc1_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_bank23_data_opc1_h.d0_0 value=0111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank23_data_opc1_h.d0_0.d = 34'b0111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_bank23_data_opc1_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank23_data_opc1_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_bank45_data_opc1_h.d0_0 value=0111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank45_data_opc1_h.d0_0.d = 34'b0111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_bank45_data_opc1_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank45_data_opc1_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_bank67_data_opc1_h.d0_0 value=0111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank67_data_opc1_h.d0_0.d = 34'b0111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_bank67_data_opc1_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_bank67_data_opc1_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_mbist0145_data_h.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_mbist0145_data_h.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_mbist0145_data_l.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_mbist0145_data_l.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_mbist2367_data_h.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_mbist2367_data_h.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdc.dff_mbist2367_data_l.d0_0 value=1111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdc.dff_mbist2367_data_l.d0_0.d = 34'b1111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq00.dff_din_hi.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq00.dff_din_hi.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq00.dff_din_lo.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq00.dff_din_lo.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq00.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq00.dff_dout.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq01.dff_din_hi.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq01.dff_din_hi.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq01.dff_din_lo.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq01.dff_din_lo.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq01.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq01.dff_dout.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq10.dff_din_hi.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq10.dff_din_hi.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq10.dff_din_lo.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq10.dff_din_lo.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq10.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq10.dff_dout.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq11.dff_din_hi.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq11.dff_din_hi.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq11.dff_din_lo.d0_0 value=111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq11.dff_din_lo.d0_0.d = 36'b111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opddq11.dff_dout.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opddq11.dff_dout.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.sio.opdhq0.dff_din_hi.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdhq0.dff_din_hi.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.sio.opdhq0.dff_din_lo.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdhq0.dff_din_lo.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.sio.opdhq1.dff_din_hi.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdhq1.dff_din_hi.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.sio.opdhq1.dff_din_lo.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opdhq1.dff_din_lo.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.sio.opds0.ff_opdhqxout.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds0.ff_opdhqxout.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds0.ff_packet_data0_h.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds0.ff_packet_data0_h.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds0.ff_packet_data0_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds0.ff_packet_data0_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds0.ff_packet_data1_h.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds0.ff_packet_data1_h.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds0.ff_packet_data1_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds0.ff_packet_data1_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds1.ff_opdhqxout.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds1.ff_opdhqxout.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds1.ff_packet_data0_h.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds1.ff_packet_data0_h.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds1.ff_packet_data0_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds1.ff_packet_data0_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds1.ff_packet_data1_h.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds1.ff_packet_data1_h.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.sio.opds1.ff_packet_data1_l.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.sio.opds1.ff_packet_data1_l.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.spc0.clk_spc.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.spc0.clk_spc.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.spc0.dec.del.exu_clkenf.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.dec.del.exu_clkenf.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.dec.del.fef.d0_0 value=0000000011111111 out=q in=d model=dff 
force tb_top.cpu.spc0.dec.del.fef.d0_0.d = 16'b0000000011111111;

// instance=tb_top.cpu.spc0.dec.del.pdisttidf.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.dec.del.pdisttidf.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.dec.del.tid_e.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.dec.del.tid_e.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.dec.del.tid_m.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.dec.del.tid_m.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.dec.del.truevalid_f.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.dec.del.truevalid_f.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.exu0.ect.fcce_ff.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.ect.fcce_ff.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.exu0.ect.fgu_tid_ff.d0_0 value=111000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.ect.fgu_tid_ff.d0_0.d = 6'b111000;

// instance=tb_top.cpu.spc0.exu0.ect.i_byp_lth.d0_0 value=1101100000000000000001100000001100000011000000110000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.ect.i_byp_lth.d0_0.d = 76'b1101100000000000000001100000001100000011000000110000000000000000000000000000;

// instance=tb_top.cpu.spc0.exu0.ect.i_estage_lth.d0_0 value=0000100000000010100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.ect.i_estage_lth.d0_0.d = 37'b0000100000000010100000000000000000000;

// instance=tb_top.cpu.spc0.exu0.ect.i_pwr0_lth.d0_0 value=10000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.ect.i_pwr0_lth.d0_0.d = 5'b10000;

// instance=tb_top.cpu.spc0.exu0.edp.i_asi0_ff.d0_0 value=10000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.edp.i_asi0_ff.d0_0.d = 65'b10000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.exu0.edp.i_misc_ff.d0_0 value=0000000000000000000000001010 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.edp.i_misc_ff.d0_0.d = 28'b0000000000000000000000001010;

// instance=tb_top.cpu.spc0.exu0.irf.i_rd_control_ff.d0_0 value=00000000000000000011 out=mq in=d model=new_dlata 
force tb_top.cpu.spc0.exu0.irf.i_rd_control_ff.d0_0.d = 20'b00000000000000000011;

// instance=tb_top.cpu.spc0.exu0.irf.i_rd_control_ff.d0_0 value=00000000000000000011 out=q in=d model=new_dlata 
force tb_top.cpu.spc0.exu0.irf.i_rd_control_ff.d0_0.d = 20'b00000000000000000011;

// instance=tb_top.cpu.spc0.exu0.irf.i_restore_ff.d0_0 value=00000000000001100 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.irf.i_restore_ff.d0_0.d = 17'b00000000000001100;

// instance=tb_top.cpu.spc0.exu0.irf.i_save_ff.d0_0 value=00000000000001100 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.irf.i_save_ff.d0_0.d = 17'b00000000000001100;

// instance=tb_top.cpu.spc0.exu0.irf.i_wr_control_ff.d0_0 value=0000000000000110 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.irf.i_wr_control_ff.d0_0.d = 16'b0000000000000110;

// instance=tb_top.cpu.spc0.exu0.rml.cansave_e2m2b2w.d0_0 value=110110110 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.cansave_e2m2b2w.d0_0.d = 9'b110110110;

// instance=tb_top.cpu.spc0.exu0.rml.cleanwin_e2m2b2w.d0_0 value=111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.cleanwin_e2m2b2w.d0_0.d = 9'b111111111;

// instance=tb_top.cpu.spc0.exu0.rml.cwp_b2w.d0_0 value=110000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.cwp_b2w.d0_0.d = 6'b110000;

// instance=tb_top.cpu.spc0.exu0.rml.cwp_m2b.d0_0 value=110000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.cwp_m2b.d0_0.d = 6'b110000;

// instance=tb_top.cpu.spc0.exu0.rml.exception_report_m2b.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.exception_report_m2b.d0_0.d = 3'b001;

// instance=tb_top.cpu.spc0.exu0.rml.i_rml_restore_en_ff.d0_0 value=000000110000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.i_rml_restore_en_ff.d0_0.d = 15'b000000110000000;

// instance=tb_top.cpu.spc0.exu0.rml.tid_p2d2e2m2b2w.d0_0 value=11111111111000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.tid_p2d2e2m2b2w.d0_0.d = 14'b11111111111000;

// instance=tb_top.cpu.spc0.exu0.rml.winblock_slot_tid_m2d2e2m.d0_0 value=111111 out=q in=d model=dff 
force tb_top.cpu.spc0.exu0.rml.winblock_slot_tid_m2d2e2m.d0_0.d = 6'b111111;

// instance=tb_top.cpu.spc0.exu1.ect.fcce_ff.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.ect.fcce_ff.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.exu1.ect.fgu_tid_ff.d0_0 value=111000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.ect.fgu_tid_ff.d0_0.d = 6'b111000;

// instance=tb_top.cpu.spc0.exu1.ect.i_byp_lth.d0_0 value=1101100000000000000001100000001100000011000000110000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.ect.i_byp_lth.d0_0.d = 76'b1101100000000000000001100000001100000011000000110000000000000000000000000000;

// instance=tb_top.cpu.spc0.exu1.ect.i_estage_lth.d0_0 value=0000100000000010100000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.ect.i_estage_lth.d0_0.d = 37'b0000100000000010100000000000000000000;

// instance=tb_top.cpu.spc0.exu1.ect.i_pwr0_lth.d0_0 value=10000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.ect.i_pwr0_lth.d0_0.d = 5'b10000;

// instance=tb_top.cpu.spc0.exu1.edp.i_asi0_ff.d0_0 value=10000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.edp.i_asi0_ff.d0_0.d = 65'b10000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.exu1.edp.i_misc_ff.d0_0 value=0000000000000000000000001010 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.edp.i_misc_ff.d0_0.d = 28'b0000000000000000000000001010;

// instance=tb_top.cpu.spc0.exu1.irf.i_rd_control_ff.d0_0 value=00000000000000000011 out=mq in=d model=new_dlata 
force tb_top.cpu.spc0.exu1.irf.i_rd_control_ff.d0_0.d = 20'b00000000000000000011;

// instance=tb_top.cpu.spc0.exu1.irf.i_rd_control_ff.d0_0 value=00000000000000000011 out=q in=d model=new_dlata 
force tb_top.cpu.spc0.exu1.irf.i_rd_control_ff.d0_0.d = 20'b00000000000000000011;

// instance=tb_top.cpu.spc0.exu1.irf.i_restore_ff.d0_0 value=00000000000001100 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.irf.i_restore_ff.d0_0.d = 17'b00000000000001100;

// instance=tb_top.cpu.spc0.exu1.irf.i_save_ff.d0_0 value=00000000000001100 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.irf.i_save_ff.d0_0.d = 17'b00000000000001100;

// instance=tb_top.cpu.spc0.exu1.irf.i_wr_control_ff.d0_0 value=0000000000000110 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.irf.i_wr_control_ff.d0_0.d = 16'b0000000000000110;

// instance=tb_top.cpu.spc0.exu1.rml.cansave_e2m2b2w.d0_0 value=110110110 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.cansave_e2m2b2w.d0_0.d = 9'b110110110;

// instance=tb_top.cpu.spc0.exu1.rml.cleanwin_e2m2b2w.d0_0 value=111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.cleanwin_e2m2b2w.d0_0.d = 9'b111111111;

// instance=tb_top.cpu.spc0.exu1.rml.cwp_b2w.d0_0 value=110000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.cwp_b2w.d0_0.d = 6'b110000;

// instance=tb_top.cpu.spc0.exu1.rml.cwp_m2b.d0_0 value=110000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.cwp_m2b.d0_0.d = 6'b110000;

// instance=tb_top.cpu.spc0.exu1.rml.exception_report_m2b.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.exception_report_m2b.d0_0.d = 3'b001;

// instance=tb_top.cpu.spc0.exu1.rml.i_rml_restore_en_ff.d0_0 value=000000110000000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.i_rml_restore_en_ff.d0_0.d = 15'b000000110000000;

// instance=tb_top.cpu.spc0.exu1.rml.tid_p2d2e2m2b2w.d0_0 value=11111111111000 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.tid_p2d2e2m2b2w.d0_0.d = 14'b11111111111000;

// instance=tb_top.cpu.spc0.exu1.rml.winblock_slot_tid_m2d2e2m.d0_0 value=111111 out=q in=d model=dff 
force tb_top.cpu.spc0.exu1.rml.winblock_slot_tid_m2d2e2m.d0_0.d = 6'b111111;

// instance=tb_top.cpu.spc0.fgu.fac.e_01.d0_0 value=0000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.e_01.d0_0.d = 37'b0000000000000000000000000000000000001;

// instance=tb_top.cpu.spc0.fgu.fac.e_02.d0_0 value=00000000111000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.e_02.d0_0.d = 17'b00000000111000000;

// instance=tb_top.cpu.spc0.fgu.fac.fb_00.d0_0 value=0000000111000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fb_00.d0_0.d = 25'b0000000111000000000000000;

// instance=tb_top.cpu.spc0.fgu.fac.fprs_frf_ctl.d0_0 value=011100000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fprs_frf_ctl.d0_0.d = 12'b011100000000;

// instance=tb_top.cpu.spc0.fgu.fac.fprs_rng.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fprs_rng.d0_0.d = 3'b100;

// instance=tb_top.cpu.spc0.fgu.fac.fw_00.d0_0 value=000111000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fw_00.d0_0.d = 21'b000111000000000000000;

// instance=tb_top.cpu.spc0.fgu.fac.fx1_00.d0_0 value=00000101100111011010000000000000000000000000000000000000000000000000000010110000000000000000000000000000000000001000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fx1_00.d0_0.d = 128'b00000101100111011010000000000000000000000000000000000000000000000000000010110000000000000000000000000000000000001000000000000000;

// instance=tb_top.cpu.spc0.fgu.fac.fx1_01.d0_0 value=000000011100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fx1_01.d0_0.d = 21'b000000011100000000000;

// instance=tb_top.cpu.spc0.fgu.fac.fx2_00.d0_0 value=0000000111000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fx2_00.d0_0.d = 16'b0000000111000000;

// instance=tb_top.cpu.spc0.fgu.fac.fx2_01.d0_0 value=000000000000000000000000000000000001000000001011000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fx2_01.d0_0.d = 60'b000000000000000000000000000000000001000000001011000000000000;

// instance=tb_top.cpu.spc0.fgu.fac.fx3_00.d0_0 value=0000000111000001000000000000100000010110000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fx3_00.d0_0.d = 52'b0000000111000001000000000000100000010110000000000000;

// instance=tb_top.cpu.spc0.fgu.fac.fx4_00.d0_0 value=0000000111000000000000100000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fx4_00.d0_0.d = 31'b0000000111000000000000100000000;

// instance=tb_top.cpu.spc0.fgu.fac.fx5_00.d0_0 value=00000001110000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.fx5_00.d0_0.d = 26'b00000001110000000000000000;

// instance=tb_top.cpu.spc0.fgu.fac.rng_6463.d0_0 value=001000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.rng_6463.d0_0.d = 6'b001000;

// instance=tb_top.cpu.spc0.fgu.fac.rng_stg1.d0_0 value=1000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fac.rng_stg1.d0_0.d = 25'b1000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fad.e_01.d0_0 value=00000000000000011100000000000000000001000010000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fad.e_01.d0_0.d = 47'b00000000000000011100000000000000000001000010000;

// instance=tb_top.cpu.spc0.fgu.fad.e_01_extra.d0_0 value=00000000000000000001100 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fad.e_01_extra.d0_0.d = 23'b00000000000000000001100;

// instance=tb_top.cpu.spc0.fgu.fdc.data_lth.d0_0 value=000000011 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdc.data_lth.d0_0.d = 9'b000000011;

// instance=tb_top.cpu.spc0.fgu.fdc.ovlf_lth.d0_0 value=0010 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdc.ovlf_lth.d0_0.d = 4'b0010;

// instance=tb_top.cpu.spc0.fgu.fdc.xrnd_lth.d0_0 value=0000011000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdc.xrnd_lth.d0_0.d = 10'b0000011000;

// instance=tb_top.cpu.spc0.fgu.fdd.ie_d00lthm1.d0_0 value=11111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdd.ie_d00lthm1.d0_0.d = 65'b11111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.fgu.fdd.ie_d00lthp1.d0_0 value=11111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdd.ie_d00lthp1.d0_0.d = 65'b11111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.fgu.fdd.ipte_clalth0.d0_0 value=00000000000000011111111100000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdd.ipte_clalth0.d0_0.d = 65'b00000000000000011111111100000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fdd.ipte_clalth1.d0_0 value=00000000000000000000000010000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdd.ipte_clalth1.d0_0.d = 65'b00000000000000000000000010000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fdd.isqe_cnt.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdd.isqe_cnt.d0_0.d = 66'b111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.fgu.fdd.isqe_flip.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fdd.isqe_flip.d0_0.d = 66'b111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.fgu.fgd.fx4_gsrtid.d0_0 value=000111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fgd.fx4_gsrtid.d0_0.d = 6'b000111;

// instance=tb_top.cpu.spc0.fgu.fic.fx2_00.d0_0 value=1100000000010000000111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fic.fx2_00.d0_0.d = 43'b1100000000010000000111111111111111111111111;

// instance=tb_top.cpu.spc0.fgu.fpc.fb_05.d0_0 value=0000000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fb_05.d0_0.d = 13'b0000000000001;

// instance=tb_top.cpu.spc0.fgu.fpc.fx1_01.d0_0 value=00111000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx1_01.d0_0.d = 8'b00111000;

// instance=tb_top.cpu.spc0.fgu.fpc.fx2_00.d0_0 value=101100110000000010000000000000000000000001010000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx2_00.d0_0.d = 51'b101100110000000010000000000000000000000001010000000;

// instance=tb_top.cpu.spc0.fgu.fpc.fx2_01.d0_0 value=10000000000010 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx2_01.d0_0.d = 14'b10000000000010;

// instance=tb_top.cpu.spc0.fgu.fpc.fx2_02.d0_0 value=00010000000001111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx2_02.d0_0.d = 17'b00010000000001111;

// instance=tb_top.cpu.spc0.fgu.fpc.fx2_05.d0_0 value=110011 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx2_05.d0_0.d = 6'b110011;

// instance=tb_top.cpu.spc0.fgu.fpc.fx3_00.d0_0 value=0010110011111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx3_00.d0_0.d = 13'b0010110011111;

// instance=tb_top.cpu.spc0.fgu.fpc.fx3_01.d0_0 value=01110000000010000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx3_01.d0_0.d = 20'b01110000000010000000;

// instance=tb_top.cpu.spc0.fgu.fpc.fx3_02.d0_0 value=0000000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx3_02.d0_0.d = 13'b0000000000001;

// instance=tb_top.cpu.spc0.fgu.fpc.fx3_03.d0_0 value=1100 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx3_03.d0_0.d = 4'b1100;

// instance=tb_top.cpu.spc0.fgu.fpc.fx3_05.d0_0 value=0000001000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx3_05.d0_0.d = 10'b0000001000;

// instance=tb_top.cpu.spc0.fgu.fpc.fx3_06.d0_0 value=0000000000000000001000001000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx3_06.d0_0.d = 28'b0000000000000000001000001000;

// instance=tb_top.cpu.spc0.fgu.fpc.fx4_00.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx4_00.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.fgu.fpc.fx4_01.d0_0 value=0000000000100000000000000000000001000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx4_01.d0_0.d = 37'b0000000000100000000000000000000001000;

// instance=tb_top.cpu.spc0.fgu.fpc.fx4_02.d0_0 value=011100000101100 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx4_02.d0_0.d = 15'b011100000101100;

// instance=tb_top.cpu.spc0.fgu.fpc.fx5_01.d0_0 value=10110001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx5_01.d0_0.d = 8'b10110001;

// instance=tb_top.cpu.spc0.fgu.fpc.fx5_02.d0_0 value=000001110000100101010000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpc.fx5_02.d0_0.d = 36'b000001110000100101010000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpe.fb_exp_res.d0_0 value=10000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpe.fb_exp_res.d0_0.d = 11'b10000000001;

// instance=tb_top.cpu.spc0.fgu.fpe.fx1_fmtsel.d0_0 value=000100100100000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpe.fx1_fmtsel.d0_0.d = 18'b000100100100000001;

// instance=tb_top.cpu.spc0.fgu.fpe.fx2_aux.d0_0 value=10000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpe.fx2_aux.d0_0.d = 11'b10000000001;

// instance=tb_top.cpu.spc0.fgu.fpe.fx2_swp_sel.d0_0 value=0000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpe.fx2_swp_sel.d0_0.d = 22'b0000000000000000000001;

// instance=tb_top.cpu.spc0.fgu.fpe.fx3_einty.d0_0 value=10000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpe.fx3_einty.d0_0.d = 11'b10000000001;

// instance=tb_top.cpu.spc0.fgu.fpe.fx4_einty.d0_0 value=001000000000110000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpe.fx4_einty.d0_0.d = 24'b001000000000110000000001;

// instance=tb_top.cpu.spc0.fgu.fpf.fb_nrd.d0_0 value=0100000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpf.fb_nrd.d0_0.d = 58'b0100000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpf.fx2_fcc.d0_0 value=01110111010010001000101010000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpf.fx2_fcc.d0_0.d = 29'b01110111010010001000101010000;

// instance=tb_top.cpu.spc0.fgu.fpf.fx3_fcc.d0_0 value=000000111000000000000010000010000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpf.fx3_fcc.d0_0.d = 54'b000000111000000000000010000010000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a0_be_ff.d0_0 value=11011111100000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a0_be_ff.d0_0.d = 41'b11011111100000000000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a0_s_ff_a.d0_0 value=1111111111111111100000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a0_s_ff_a.d0_0.d = 40'b1111111111111111100000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a10_x_ff_a.d0_0 value=01111001111111111111111000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a10_x_ff_a.d0_0.d = 44'b01111001111111111111111000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a1_be_ff.d0_0 value=1111111111000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a1_be_ff.d0_0.d = 64'b1111111111000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a1_s_ff_a.d0_0 value=11111111111111111100000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a1_s_ff_a.d0_0.d = 41'b11111111111111111100000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a2_be_ff_a.d0_0 value=1111111111111111111110000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a2_be_ff_a.d0_0.d = 31'b1111111111111111111110000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a2_s_ff_a.d0_0 value=11111111111111111100000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a2_s_ff_a.d0_0.d = 41'b11111111111111111100000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a32_x_ff_a.d0_0 value=11111001111111111111000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a32_x_ff_a.d0_0.d = 44'b11111001111111111111000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a3_be_ff.d0_0 value=111111111100000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a3_be_ff.d0_0.d = 63'b111111111100000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a3_c_ff_a.d0_0 value=0000000000000100000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a3_c_ff_a.d0_0.d = 37'b0000000000000100000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a3_s_ff_a.d0_0 value=111111111111110000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a3_s_ff_a.d0_0.d = 39'b111111111111110000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a4_c_hi_ff.d0_0 value=000000000000000000000000000000000000000000000000000000000001000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a4_c_hi_ff.d0_0.d = 69'b000000000000000000000000000000000000000000000000000000000001000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_a4_s_hi_ff.d0_0 value=111111111111111111111111111111111111111111111111111111111111111000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_a4_s_hi_ff.d0_0.d = 72'b111111111111111111111111111111111111111111111111111111111111111000000000;

// instance=tb_top.cpu.spc0.fgu.fpy.i_fx5_ff.d0_0 value=11000000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.fpy.i_fx5_ff.d0_0.d = 68'b11000000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.fgu.frf.frf_read_ctl_in2ph2.d0_0 value=000000000000111 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.frf.frf_read_ctl_in2ph2.d0_0.d = 15'b000000000000111;

// instance=tb_top.cpu.spc0.fgu.frf.frf_write_input_ctl_in2fb.d0_0 value=11100000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.fgu.frf.frf_write_input_ctl_in2fb.d0_0.d = 20'b11100000000000000000;

// instance=tb_top.cpu.spc0.gkt.ipc.dff_ncu_pb.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipc.dff_ncu_pb.d0_0.d = 5'b01111;

// instance=tb_top.cpu.spc0.gkt.ipc.dff_pb_sel.d0_0 value=100100 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipc.dff_pb_sel.d0_0.d = 6'b100100;

// instance=tb_top.cpu.spc0.gkt.ipc.dff_req_drop_latx.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipc.dff_req_drop_latx.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.gkt.ipc.dff_unit_ndrop_pa.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipc.dff_unit_ndrop_pa.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.gkt.ipd.i_ifu_addr_v0_muxreg.d0_0 value=010000100000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipd.i_ifu_addr_v0_muxreg.d0_0.d = 66'b010000100000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.gkt.ipd.i_mmu_addr_v0_muxreg.d0_0 value=001000100000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipd.i_mmu_addr_v0_muxreg.d0_0.d = 66'b001000100000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.gkt.ipd.i_ncu_reg.d0_0 value=001111 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipd.i_ncu_reg.d0_0.d = 6'b001111;

// instance=tb_top.cpu.spc0.gkt.ipd.i_req_li_reg.d0_0 value=1000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipd.i_req_li_reg.d0_0.d = 19'b1000000000000000000;

// instance=tb_top.cpu.spc0.gkt.ipd.i_spu_addr_v0_muxreg.d0_0 value=000100100000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.gkt.ipd.i_spu_addr_v0_muxreg.d0_0.d = 66'b000100100000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.ifu_cmu.lsc.lsc_cpkt_reg.d0_0 value=00000010000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_cmu.lsc.lsc_cpkt_reg.d0_0.d = 11'b00000010000;

// instance=tb_top.cpu.spc0.ifu_cmu.lsd.paddr_lat.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_cmu.lsd.paddr_lat.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.any_instr_v_c_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.any_instr_v_c_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.br_misp_data_dup_reg.d0_0 value=111111110000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.br_misp_data_dup_reg.d0_0.d = 12'b111111110000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.br_misp_data_reg.d0_0 value=11110000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.br_misp_data_reg.d0_0.d = 8'b11110000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.bus_first_reg.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.bus_first_reg.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.ic_instr_v_reg.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.ic_instr_v_reg.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.inv_way1_bf_reg.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.inv_way1_bf_reg.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.inv_way_bf_reg.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.inv_way_bf_reg.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_1_reg.d0_0 value=10000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_1_reg.d0_0.d = 5'b10000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_2_reg.d0_0 value=10000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_2_reg.d0_0.d = 5'b10000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_in_reg.d0_0 value=10000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_in_reg.d0_0.d = 5'b10000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.mbist_output.d0_0 value=100100 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.mbist_output.d0_0.d = 6'b100100;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr0_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr0_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr1_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr1_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr2_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr2_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr3_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr3_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr4_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr4_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr5_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr5_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr6_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr6_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr7_pc_f_inc_reg.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr7_pc_f_inc_reg.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr_c_ic_disable_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr_c_ic_disable_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.tid_dec_w_reg.d0_0 value=10001000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.tid_dec_w_reg.d0_0.d = 8'b10001000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.wrway_bf_reg.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.wrway_bf_reg.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_asi_ctl.rng_stg2_ctl.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_asi_ctl.rng_stg2_ctl.d0_0.d = 3'b100;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_asi_ctl.rng_stg2_decctl.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_asi_ctl.rng_stg2_decctl.d0_0.d = 2'b10;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_byp_dp.itb_data_for_cam.d0_0 value=0000000000000010 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_byp_dp.itb_data_for_cam.d0_0.d = 16'b0000000000000010;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_cms_ctl.rep_way_reg.d0_0 value=0000000100 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_cms_ctl.rep_way_reg.d0_0.d = 10'b0000000100;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.br_tid_reg.d0_0 value=111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.br_tid_reg.d0_0.d = 12'b111111111111;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.itlb_probe_l_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.itlb_probe_l_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.pstate_am_reg.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.pstate_am_reg.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.tid_dec_w_reg.d0_0 value=10001000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.tid_dec_w_reg.d0_0.d = 8'b10001000;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.index_reg_i.d0_0 value=111111111 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.index_reg_i.d0_0.d = 9'b111111111;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.quad_en_reg.d0_0 value=0000 out=q_l in=d model=msffi 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.quad_en_reg.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.rdreq_reg.d0_0 value=1 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.rdreq_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.way_c_reg.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.way_c_reg.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.way_f_reg.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.way_f_reg.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrreq_reg.d0_0 value=1 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrreq_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_0_reg.d0_0 value=1 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_0_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_1_reg.d0_0 value=1 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_1_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_2_reg.d0_0 value=1 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_2_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.cache_way_hit_reg.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.cache_way_hit_reg.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tlb_cam_hit_reg.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tlb_cam_hit_reg.d0_0.d = 3'b100;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tte_tag_out_reg.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tte_tag_out_reg.d0_0.d = 66'b111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tte_u_bit_out_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tte_u_bit_out_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_itc_ctl.itc_sel_demap_reg.d0_0 value=0000010 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_itc_ctl.itc_sel_demap_reg.d0_0.d = 7'b0000010;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_itc_ctl.tte1_lat.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_itc_ctl.tte1_lat.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_itd_dp.tte1_lat.d0_0 value=00000000000000000000000000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_itd_dp.tte1_lat.d0_0.d = 59'b00000000000000000000000000000000000000000000000000000000001;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm0.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm0.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm1.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm1.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm2.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm2.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm3.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm3.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm4.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm4.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm5.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm5.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm6.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm6.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm7.ignore_by_pass_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm7.ignore_by_pass_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ftu.hdr.sram_header_instance.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ftu.hdr.sram_header_instance.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq0.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq0.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq0.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq0.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq1.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq1.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq1.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq1.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq2.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq2.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq2.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq2.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq3.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq3.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq3.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq3.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq4.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq4.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq4.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq4.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq5.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq5.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq5.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq5.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq6.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq6.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq6.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq6.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq7.buff_clken_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq7.buff_clken_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.ifu_ibu.ibq7.fetch_sig_reg.d0_0 value=00100000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.ifu_ibu.ibq7.fetch_sig_reg.d0_0.d = 14'b00100000000000;

// instance=tb_top.cpu.spc0.lsu.ard.i_rngl_stg1_reg.d0_0 value=10000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.ard.i_rngl_stg1_reg.d0_0.d = 65'b10000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.lsu.asc.ascl_vld_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.asc.ascl_vld_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.lsu.asc.hole_count.d0_0 value=1001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.asc.hole_count.d0_0.d = 4'b1001;

// instance=tb_top.cpu.spc0.lsu.cic.dff_cpq_sel.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.cic.dff_cpq_sel.d0_0.d = 2'b10;

// instance=tb_top.cpu.spc0.lsu.dac.dff_baddr_b.d0_0 value=0000000101 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dac.dff_baddr_b.d0_0.d = 10'b0000000101;

// instance=tb_top.cpu.spc0.lsu.dac.dff_endian_b.d0_0 value=01 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dac.dff_endian_b.d0_0.d = 2'b01;

// instance=tb_top.cpu.spc0.lsu.dac.dff_ld_sz_b.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dac.dff_ld_sz_b.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.lsu.dca.dff_ctl_b.d0_0 value=10001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dca.dff_ctl_b.d0_0.d = 5'b10001;

// instance=tb_top.cpu.spc0.lsu.dca.dff_ctl_m_1.d0_0 value=1111111111111111 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.lsu.dca.dff_ctl_m_1.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.spc0.lsu.dca.lat_ctl_eb.d0_0 value=0000001 out=latout in=d model=tisram_msff 
force tb_top.cpu.spc0.lsu.dca.lat_ctl_eb.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_asi_b.d0_0 value=000000100000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_asi_b.d0_0.d = 24'b000000100000000000000000;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_asi_m.d0_0 value=000100000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_asi_m.d0_0.d = 12'b000100000000;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_excp_b.d0_0 value=00011 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_excp_b.d0_0.d = 5'b00011;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_new_lru_w.d0_0 value=0001110000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_new_lru_w.d0_0.d = 13'b0001110000000;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_pwr_mgmt.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_pwr_mgmt.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_sba_par.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_sba_par.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_tid_b.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_tid_b.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_tid_e.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_tid_e.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_tid_m.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_tid_m.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.lsu.dcc.dff_tid_w.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcc.dff_tid_w.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.lsu.dcs.dff_context_m.d0_0 value=10000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dcs.dff_context_m.d0_0.d = 14'b10000000000000;

// instance=tb_top.cpu.spc0.lsu.dva.dff_din.d0_0 value=11111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.dva.dff_din.d0_0.d = 32'b11111111111111111111111111111111;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_inst_b.d0_0 value=000111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_inst_b.d0_0.d = 6'b000111;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_ld_inst_e.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_ld_inst_e.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_ld_lmq_en_b.d0_0 value=001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_ld_lmq_en_b.d0_0.d = 3'b001;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w.d0_0 value=0111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w.d0_0.d = 4'b0111;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w2.d0_0 value=0111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w2.d0_0.d = 4'b0111;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w3.d0_0 value=0111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w3.d0_0.d = 4'b0111;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_ld_sel.d0_0 value=1000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_ld_sel.d0_0.d = 10'b1000000000;

// instance=tb_top.cpu.spc0.lsu.lmc.dff_thread_w.d0_0 value=10000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lmc.dff_thread_w.d0_0.d = 8'b10000000;

// instance=tb_top.cpu.spc0.lsu.lru.dff_bit_en.d0_0 value=00000000000000000000000011111111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lru.dff_bit_en.d0_0.d = 32'b00000000000000000000000011111111;

// instance=tb_top.cpu.spc0.lsu.lru.dff_din.d0_0 value=00000111000001110000011100000111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.lru.dff_din.d0_0.d = 32'b00000111000001110000011100000111;

// instance=tb_top.cpu.spc0.lsu.pic.dff_asi_pm.d0_0 value=100000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.pic.dff_asi_pm.d0_0.d = 6'b100000;

// instance=tb_top.cpu.spc0.lsu.pic.dff_asi_req.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.pic.dff_asi_req.d0_0.d = 3'b010;

// instance=tb_top.cpu.spc0.lsu.red.sram_header_instance.ff_io_cmp_sync_en.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.red.sram_header_instance.ff_io_cmp_sync_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.lsu.sbc.dff_cam_hit.d0_0 value=111000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbc.dff_cam_hit.d0_0.d = 9'b111000000;

// instance=tb_top.cpu.spc0.lsu.sbc.dff_stb_err.d0_0 value=0000000110 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbc.dff_stb_err.d0_0.d = 10'b0000000110;

// instance=tb_top.cpu.spc0.lsu.sbc.dff_thread_b.d0_0 value=10000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbc.dff_thread_b.d0_0.d = 8'b10000000;

// instance=tb_top.cpu.spc0.lsu.sbc.dff_tid_m.d0_0 value=111111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbc.dff_tid_m.d0_0.d = 6'b111111;

// instance=tb_top.cpu.spc0.lsu.sbs0.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs0.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sbs1.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs1.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sbs2.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs2.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sbs3.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs3.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sbs4.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs4.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sbs5.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs5.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sbs6.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs6.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sbs7.dff_asi_pipe.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sbs7.dff_asi_pipe.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.lsu.sec.dff_cparity.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sec.dff_cparity.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.lsu.sec.dff_st_sz.d0_0 value=00000000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sec.dff_st_sz.d0_0.d = 14'b00000000000001;

// instance=tb_top.cpu.spc0.lsu.sed.dff_prty_bits.d0_0 value=11101111000011000100000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sed.dff_prty_bits.d0_0.d = 26'b11101111000011000100000000;

// instance=tb_top.cpu.spc0.lsu.sed.dff_rd_data_0.d0_0 value=111111111111111111111111101111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sed.dff_rd_data_0.d0_0.d = 42'b111111111111111111111111101111111111111111;

// instance=tb_top.cpu.spc0.lsu.sed.dff_rd_data_1.d0_0 value=111111111111111111111111101111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.sed.dff_rd_data_1.d0_0.d = 42'b111111111111111111111111101111111111111111;

// instance=tb_top.cpu.spc0.lsu.stb_cam.cam_tid_din.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.stb_cam.cam_tid_din.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.lsu.stb_cam.camwr_din.d0_0 value=0000000000000000000000000000000000000100000000 out=latout in=d model=scm_msff_lat 
force tb_top.cpu.spc0.lsu.stb_cam.camwr_din.d0_0.d = 46'b0000000000000000000000000000000000000100000000;

// instance=tb_top.cpu.spc0.lsu.stb_cam.camwr_din.d0_0 value=0000000000000000000000000000000000000100000000 out=q in=d model=scm_msff_lat 
force tb_top.cpu.spc0.lsu.stb_cam.camwr_din.d0_0.d = 46'b0000000000000000000000000000000000000100000000;

// instance=tb_top.cpu.spc0.lsu.stb_ram.dff_din_lo.d0_0 value=000000000000000000000000000000000000000001 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.stb_ram.dff_din_lo.d0_0.d = 42'b000000000000000000000000000000000000000001;

// instance=tb_top.cpu.spc0.lsu.stb_ram.dff_wr_addr.d0_0 value=111000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.stb_ram.dff_wr_addr.d0_0.d = 6'b111000;

// instance=tb_top.cpu.spc0.lsu.tgd.dff_va_b.d0_0 value=000000000000000000000000000000000000000000000111100 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tgd.dff_va_b.d0_0.d = 51'b000000000000000000000000000000000000000000000111100;

// instance=tb_top.cpu.spc0.lsu.tlb.cache_way_hit_reg.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlb.cache_way_hit_reg.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.lsu.tlb.cam_ctl_lat.d0_0 value=00000000000000001000000000000000000000000000000000000000000000000010000000 out=mq in=d model=new_dlata 
force tb_top.cpu.spc0.lsu.tlb.cam_ctl_lat.d0_0.d = 74'b00000000000000001000000000000000000000000000000000000000000000000010000000;

// instance=tb_top.cpu.spc0.lsu.tlb.cam_ctl_lat.d0_0 value=00000000000000001000000000000000000000000000000000000000000000000010000000 out=q in=d model=new_dlata 
force tb_top.cpu.spc0.lsu.tlb.cam_ctl_lat.d0_0.d = 74'b00000000000000001000000000000000000000000000000000000000000000000010000000;

// instance=tb_top.cpu.spc0.lsu.tlb.pa_reg.d0_0 value=111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlb.pa_reg.d0_0.d = 27'b111111111111111111111111111;

// instance=tb_top.cpu.spc0.lsu.tlb.page_size_mask_reg.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlb.page_size_mask_reg.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.lsu.tlb.tlb_cam_hit_reg.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlb.tlb_cam_hit_reg.d0_0.d = 3'b100;

// instance=tb_top.cpu.spc0.lsu.tlb.tte_data_reg.d0_0 value=10000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlb.tte_data_reg.d0_0.d = 38'b10000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.lsu.tlb.tte_tag_out_reg.d0_0 value=111111111111111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlb.tte_tag_out_reg.d0_0.d = 66'b111111111111111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.lsu.tlb.tte_u_bit_out_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlb.tte_u_bit_out_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.lsu.tlc.wr_vld_latch.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tlc.wr_vld_latch.d0_0.d = 3'b010;

// instance=tb_top.cpu.spc0.lsu.tld.tte2_lat.d0_0 value=0001000000000000010000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.lsu.tld.tte2_lat.d0_0.d = 52'b0001000000000000010000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mb0.cntl_reg.d0_0 value=0100000001111111000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mb0.cntl_reg.d0_0.d = 28'b0100000001111111000000000000;

// instance=tb_top.cpu.spc0.mb0.exp_stb_cam_hit_delay.d0_0 value=111 out=q in=d model=dff 
force tb_top.cpu.spc0.mb0.exp_stb_cam_hit_delay.d0_0.d = 3'b111;

// instance=tb_top.cpu.spc0.mb0.input_signals_reg.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.spc0.mb0.input_signals_reg.d0_0.d = 2'b10;

// instance=tb_top.cpu.spc0.mb0.pmen.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.spc0.mb0.pmen.d0_0.d = 3'b010;

// instance=tb_top.cpu.spc0.mb1.cntl_reg.d0_0 value=010000000111111100000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mb1.cntl_reg.d0_0.d = 24'b010000000111111100000000;

// instance=tb_top.cpu.spc0.mb1.input_signals_reg.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.spc0.mb1.input_signals_reg.d0_0.d = 2'b10;

// instance=tb_top.cpu.spc0.mb1.out_cmp_sel_reg.d0_0 value=00001 out=q in=d model=dff 
force tb_top.cpu.spc0.mb1.out_cmp_sel_reg.d0_0.d = 5'b00001;

// instance=tb_top.cpu.spc0.mb1.pmen.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.spc0.mb1.pmen.d0_0.d = 3'b010;

// instance=tb_top.cpu.spc0.mb2.cntl_reg.d0_0 value=01000011111111110000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mb2.cntl_reg.d0_0.d = 29'b01000011111111110000000000000;

// instance=tb_top.cpu.spc0.mb2.input_signals_reg.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.spc0.mb2.input_signals_reg.d0_0.d = 2'b10;

// instance=tb_top.cpu.spc0.mb2.pmen.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.spc0.mb2.pmen.d0_0.d = 3'b010;

// instance=tb_top.cpu.spc0.mmu.ase.lsu_context_w_lat.d0_0 value=0000000001000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.ase.lsu_context_w_lat.d0_0.d = 25'b0000000001000000000000000;

// instance=tb_top.cpu.spc0.mmu.asi.mbist_cmpsel_2_lat.d0_0 value=01 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.mbist_cmpsel_2_lat.d0_0.d = 2'b01;

// instance=tb_top.cpu.spc0.mmu.asi.mbist_cmpsel_lat.d0_0 value=01 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.mbist_cmpsel_lat.d0_0.d = 2'b01;

// instance=tb_top.cpu.spc0.mmu.asi.rd_tte_lat.d0_0 value=0000000000000000100000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.rd_tte_lat.d0_0.d = 25'b0000000000000000100000000;

// instance=tb_top.cpu.spc0.mmu.asi.stg1_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.stg1_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.mmu.asi.stg2_ctl_lat.d0_0 value=1000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.stg2_ctl_lat.d0_0.d = 16'b1000000000000000;

// instance=tb_top.cpu.spc0.mmu.asi.stg2_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.stg2_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.mmu.asi.stg3_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.stg3_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.mmu.asi.stg4_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.stg4_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.mmu.asi.tag_access_tid_0_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.tag_access_tid_0_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.mmu.asi.tag_access_tid_1_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.asi.tag_access_tid_1_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.mmu.htc.gkt_hw0_lat0.d0_0 value=0000000000001000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.gkt_hw0_lat0.d0_0.d = 19'b0000000000001000000;

// instance=tb_top.cpu.spc0.mmu.htc.hw4_stg_lat1.d0_0 value=00100000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.hw4_stg_lat1.d0_0.d = 8'b00100000;

// instance=tb_top.cpu.spc0.mmu.htc.hw4_stg_lat2.d0_0 value=1111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.hw4_stg_lat2.d0_0.d = 16'b1111111111111111;

// instance=tb_top.cpu.spc0.mmu.htc.m1_stg_lat.d0_0 value=000010 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.m1_stg_lat.d0_0.d = 6'b000010;

// instance=tb_top.cpu.spc0.mmu.htc.m2_stg_lat2.d0_0 value=00000001000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.m2_stg_lat2.d0_0.d = 17'b00000001000000000;

// instance=tb_top.cpu.spc0.mmu.htc.m3_stg_lat1.d0_0 value=0000000000010 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.m3_stg_lat1.d0_0.d = 13'b0000000000010;

// instance=tb_top.cpu.spc0.mmu.htc.rr_addr_hw2_lat.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.rr_addr_hw2_lat.d0_0.d = 3'b100;

// instance=tb_top.cpu.spc0.mmu.htc.stg_hw3_lat.d0_0 value=00100 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htc.stg_hw3_lat.d0_0.d = 5'b00100;

// instance=tb_top.cpu.spc0.mmu.htd.e0_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e0_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.e1_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e1_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.e2_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e2_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.e3_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e3_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.e4_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e4_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.e5_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e5_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.e6_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e6_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.e7_tte_reg_w40.d0_0 value=1000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.e7_tte_reg_w40.d0_0.d = 40'b1000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.mmu.htd.reg_offsethw4_w27.d0_0 value=111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.reg_offsethw4_w27.d0_0.d = 27'b111111111111111111111111111;

// instance=tb_top.cpu.spc0.mmu.htd.reg_rangehw4_w55.d0_0 value=1111111111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.reg_rangehw4_w55.d0_0.d = 55'b1111111111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.mmu.htd.reg_tsbconf_m2_w39.d0_0 value=111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.htd.reg_tsbconf_m2_w39.d0_0.d = 39'b111111111111111111111111111111111111111;

// instance=tb_top.cpu.spc0.mmu.mel0.ecc_lat.d0_0 value=1100 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.mel0.ecc_lat.d0_0.d = 4'b1100;

// instance=tb_top.cpu.spc0.mmu.mel1.ecc_lat.d0_0 value=1100 out=q in=d model=dff 
force tb_top.cpu.spc0.mmu.mel1.ecc_lat.d0_0.d = 4'b1100;

// instance=tb_top.cpu.spc0.msf0.bank2_lat.d0_0 value=100 out=q in=d model=dff 
force tb_top.cpu.spc0.msf0.bank2_lat.d0_0.d = 3'b100;

// instance=tb_top.cpu.spc0.msf0.bank4_lat.d0_0 value=0010 out=q in=d model=dff 
force tb_top.cpu.spc0.msf0.bank4_lat.d0_0.d = 4'b0010;

// instance=tb_top.cpu.spc0.pku.swl0.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl0.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl0.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl0.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl0.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl0.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl1.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl1.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl1.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl1.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl1.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl1.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl2.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl2.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl2.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl2.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl2.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl2.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl3.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl3.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl3.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl3.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl3.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl3.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl4.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl4.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl4.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl4.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl4.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl4.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl5.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl5.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl5.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl5.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl5.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl5.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl6.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl6.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl6.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl6.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl6.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl6.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl7.not_annul_ds1_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl7.not_annul_ds1_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl7.not_annul_ds2_f.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl7.not_annul_ds2_f.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pku.swl7.readyf.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.pku.swl7.readyf.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.pmu.pmu_pct_ctl.asi.d0_0 value=00000000000110 out=q in=d model=dff 
force tb_top.cpu.spc0.pmu.pmu_pct_ctl.asi.d0_0.d = 14'b00000000000110;

// instance=tb_top.cpu.spc0.pmu.pmu_pct_ctl.events.d0_0 value=011000010000001100001000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.pmu.pmu_pct_ctl.events.d0_0.d = 66'b011000010000001100001000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.pmu.pmu_pct_ctl.lsu_e2m.d0_0 value=0000000000000000000001000100 out=q in=d model=dff 
force tb_top.cpu.spc0.pmu.pmu_pct_ctl.lsu_e2m.d0_0.d = 28'b0000000000000000000001000100;

// instance=tb_top.cpu.spc0.pmu.pmu_pct_ctl.lsutid.d0_0 value=100100100 out=q in=d model=dff 
force tb_top.cpu.spc0.pmu.pmu_pct_ctl.lsutid.d0_0.d = 9'b100100100;

// instance=tb_top.cpu.spc0.pmu.pmu_pct_ctl.pic_st.d0_0 value=00000101 out=q in=d model=dff 
force tb_top.cpu.spc0.pmu.pmu_pct_ctl.pic_st.d0_0.d = 8'b00000101;

// instance=tb_top.cpu.spc0.pmu.pmu_pct_ctl.pwrm.d0_0 value=00100 out=q in=d model=dff 
force tb_top.cpu.spc0.pmu.pmu_pct_ctl.pwrm.d0_0.d = 5'b00100;

// instance=tb_top.cpu.spc0.tlu.asi.compare_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.compare_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.asi.mbist_cmpsel_2_lat.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.mbist_cmpsel_2_lat.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.tlu.asi.mbist_cmpsel_lat.d0_0 value=0001 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.mbist_cmpsel_lat.d0_0.d = 4'b0001;

// instance=tb_top.cpu.spc0.tlu.asi.rng_stg4.d0_0 value=10000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.rng_stg4.d0_0.d = 65'b10000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.tlu.asi.stg1_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.stg1_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.asi.stg2_ctl_lat.d0_0 value=100000000000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.stg2_ctl_lat.d0_0.d = 72'b100000000000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.tlu.asi.stg2_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.stg2_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.asi.stg3_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.stg3_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.asi.stg4_en_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.stg4_en_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.asi.wr_tid_dec_lat.d0_0 value=00000001 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.asi.wr_tid_dec_lat.d0_0.d = 8'b00000001;

// instance=tb_top.cpu.spc0.tlu.cep.asi_lat.d0_0 value=1000000000000000000000000000000000000000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.cep.asi_lat.d0_0.d = 64'b1000000000000000000000000000000000000000000000000000000000000000;

// instance=tb_top.cpu.spc0.tlu.fls0.fast_tid_dec_b_lat.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls0.fast_tid_dec_b_lat.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.tlu.fls0.hpriv_bar_or_ie_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls0.hpriv_bar_or_ie_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.fls0.l1en_b2w_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls0.l1en_b2w_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.fls0.l_real_w_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls0.l_real_w_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.fls0.tid_b_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls0.tid_b_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.fls0.tl_eq_0_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls0.tl_eq_0_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.fls1.fast_tid_dec_b_lat.d0_0 value=1000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls1.fast_tid_dec_b_lat.d0_0.d = 4'b1000;

// instance=tb_top.cpu.spc0.tlu.fls1.hpriv_bar_or_ie_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls1.hpriv_bar_or_ie_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.fls1.l1en_b2w_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls1.l1en_b2w_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.fls1.l_real_w_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls1.l_real_w_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.fls1.tid_b_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls1.tid_b_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.fls1.tl_eq_0_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.fls1.tl_eq_0_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.ras.s_dsfar_lat.d0_0 value=11000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.ras.s_dsfar_lat.d0_0.d = 5'b11000;

// instance=tb_top.cpu.spc0.tlu.ras.tid0_b_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.ras.tid0_b_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.ras.tid0_w1_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.ras.tid0_w1_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.ras.tid0_w_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.ras.tid0_w_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.ras.tid1_b_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.ras.tid1_b_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.ras.tid1_w1_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.ras.tid1_w1_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.ras.tid1_w_lat.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.ras.tid1_w_lat.d0_0.d = 2'b11;

// instance=tb_top.cpu.spc0.tlu.tca.dff_din_hi.d0_0 value=110001111000000000000000000000000000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.tca.dff_din_hi.d0_0.d = 36'b110001111000000000000000000000000000;

// instance=tb_top.cpu.spc0.tlu.tca.dff_rd_en.d0_0 value=1 out=mq in=d model=new_dlata 
force tb_top.cpu.spc0.tlu.tca.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.tca.dff_rd_en.d0_0 value=1 out=q in=d model=new_dlata 
force tb_top.cpu.spc0.tlu.tca.dff_rd_en.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.tel0.ecc_lat.d0_0 value=11111111111111110000000111111101111111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.tel0.ecc_lat.d0_0.d = 38'b11111111111111110000000111111101111111;

// instance=tb_top.cpu.spc0.tlu.tel1.ecc_lat.d0_0 value=11111111111111110000000111111101111111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.tel1.ecc_lat.d0_0.d = 38'b11111111111111110000000111111101111111;

// instance=tb_top.cpu.spc0.tlu.trl0.gl_rest_lat.d0_0 value=1110 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl0.gl_rest_lat.d0_0.d = 4'b1110;

// instance=tb_top.cpu.spc0.tlu.trl0.l1en_per_thread_int_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl0.l1en_per_thread_int_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.trl0.p_quiesce_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl0.p_quiesce_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.trl0.pre_allow_don_ret_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl0.pre_allow_don_ret_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.trl0.pre_allow_trap_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl0.pre_allow_trap_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.trl0.stb_empty_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl0.stb_empty_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.trl0.tic_compare_lat.d0_0 value=100000 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl0.tic_compare_lat.d0_0.d = 6'b100000;

// instance=tb_top.cpu.spc0.tlu.trl1.gl_rest_lat.d0_0 value=1110 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl1.gl_rest_lat.d0_0.d = 4'b1110;

// instance=tb_top.cpu.spc0.tlu.trl1.l1en_per_thread_int_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl1.l1en_per_thread_int_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.trl1.p_quiesce_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl1.p_quiesce_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.spc0.tlu.trl1.pre_allow_don_ret_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl1.pre_allow_don_ret_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.trl1.pre_allow_trap_lat.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl1.pre_allow_trap_lat.d0_0.d = 1'b1;

// instance=tb_top.cpu.spc0.tlu.trl1.stb_empty_lat.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.spc0.tlu.trl1.stb_empty_lat.d0_0.d = 4'b1111;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.alatch value=1 out=q in=d model=cl_sc1_alatch_4x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.alatch.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.blatch_divr value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.blatch_divr.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.ccu_div_ph_flop value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.ccu_div_ph_flop.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.observe_flops.obs_ff2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.observe_flops.obs_ff2.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.clk_stopper.blatch value=1 out=latout in=d model=cl_sc1_blatch_4x 
force tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.clk_stopper.blatch.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.por_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.por_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.por_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.por_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg1 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d = 1'b1;

// instance=tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg2 value=1 out=q in=d model=cl_sc1_msff_1x 
force tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_bnkstop_reg.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_bnkstop_reg.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_cmpsync_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_cmpsync_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_l2tstop_reg.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_l2tstop_reg.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_mcudrstop_reg.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_mcudrstop_reg.d0_0.d = 4'b1111;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_mcufbdstop_reg.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_mcufbdstop_reg.d0_0.d = 4'b1111;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_mcuiostop_reg.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_mcuiostop_reg.d0_0.d = 4'b1111;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_mcustop_reg.d0_0 value=1111 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_mcustop_reg.d0_0.d = 4'b1111;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_soc0iostop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_soc0iostop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_soc0stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_soc0stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_soc1iostop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_soc1iostop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_soc2iostop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_soc2iostop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_soc3iostop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_soc3iostop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_soc3stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_soc3stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc0stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc0stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc1stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc1stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc2stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc2stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc3stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc3stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc4stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc4stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc5stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc5stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc6stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc6stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.clkstp_ctl.clkstp_spc7stop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.clkstp_ctl.clkstp_spc7stop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.mbist_ctl.bank_avail_reg.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.bank_avail_reg.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.tcu.mbist_ctl.bank_enable_status_reg.d0_0 value=01111 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.bank_enable_status_reg.d0_0.d = 5'b01111;

// instance=tb_top.cpu.tcu.mbist_ctl.core_avail_reg.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.core_avail_reg.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.tcu.mbist_ctl.core_enable_status_reg.d0_0 value=11111111 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.core_enable_status_reg.d0_0.d = 8'b11111111;

// instance=tb_top.cpu.tcu.mbist_ctl.csr_mbist_mode_reg.d0_0 value=0010 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.csr_mbist_mode_reg.d0_0.d = 4'b0010;

// instance=tb_top.cpu.tcu.mbist_ctl.csr_ucb_data_reg.d0_0 value=0000000000000000000000000000000000000000000000000000000000000010 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.csr_ucb_data_reg.d0_0.d = 64'b0000000000000000000000000000000000000000000000000000000000000010;

// instance=tb_top.cpu.tcu.mbist_ctl.dmo_ctl.dmo_dmodf_reg.d0_0 value=010 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.dmo_ctl.dmo_dmodf_reg.d0_0.d = 3'b010;

// instance=tb_top.cpu.tcu.mbist_ctl.mbist_done_fail_reg.d0_0 value=10 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.mbist_done_fail_reg.d0_0.d = 2'b10;

// instance=tb_top.cpu.tcu.mbist_ctl.mbist_done_reg.d0_0 value=111111111111111111111111111111111111111111111111 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.mbist_done_reg.d0_0.d = 48'b111111111111111111111111111111111111111111111111;

// instance=tb_top.cpu.tcu.mbist_ctl.tcu_mbist_sync_en_reg.d0_0 value=101 out=q in=d model=dff 
force tb_top.cpu.tcu.mbist_ctl.tcu_mbist_sync_en_reg.d0_0.d = 3'b101;

// instance=tb_top.cpu.tcu.regs_ctl.spare_flops.d0_0 value=000010000 out=q in=d model=dff 
force tb_top.cpu.tcu.regs_ctl.spare_flops.d0_0.d = 9'b000010000;

// instance=tb_top.cpu.tcu.regs_ctl.tcuregs_cmpiosync_reg.d0_0 value=101 out=q in=d model=dff 
force tb_top.cpu.tcu.regs_ctl.tcuregs_cmpiosync_reg.d0_0.d = 3'b101;

// instance=tb_top.cpu.tcu.regs_ctl.tcuregs_ttstart_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.regs_ctl.tcuregs_ttstart_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk0_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk0_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk1_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk1_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk2_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk2_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk3_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk3_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk4_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk4_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk5_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk5_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk6_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk6_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk7_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk7_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu0_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu0_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu1_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu1_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu2_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu2_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu3_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu3_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc0_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc0_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc1_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc1_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc2_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc2_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc3_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc3_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc0_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc0_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc1_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc1_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc2_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc2_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc3_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc3_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc4_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc4_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc5_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc5_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc6_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc6_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc7_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc7_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk0_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk0_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk1_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk1_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk1_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk1_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk2_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk2_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk2_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk2_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk3_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk3_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk4_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk4_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk4_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk4_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk5_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk5_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk5_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk5_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk6_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk6_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk6_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk6_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk7_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk7_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk7_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk7_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t0_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t0_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t1_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t1_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t1_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t1_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t2_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t2_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t2_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t2_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t3_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t3_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t4_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t4_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t4_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t4_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t5_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t5_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t5_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t5_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t6_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t6_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t6_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t6_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t7_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t7_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t7_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t7_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu0_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu0_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu1_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu1_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu1_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu1_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu2_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu2_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu2_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu2_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu3_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu3_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc0_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc0_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc1_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc1_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc2_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc2_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc3_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc3_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc0_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc0_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc1_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc1_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc1_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc1_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc2_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc2_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc2_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc2_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc3_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc3_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc4_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc4_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc4_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc4_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc5_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc5_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc5_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc5_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc6_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc6_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc6_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc6_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc7_0.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc7_0.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc7_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc7_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu1_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu1_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu2_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu2_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu1_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu1_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu2_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu2_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc0_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc0_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc1_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc1_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc2_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc2_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc3_1.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc3_1.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_cesq_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_cesq_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_cmpdrsync_reg.d0_0 value=011 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_cmpdrsync_reg.d0_0.d = 3'b011;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_cntdly_reg.d0_0 value=1111100 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_cntdly_reg.d0_0.d = 7'b1111100;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_cntstart_reg.d0_0 value=0000001 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_cntstart_reg.d0_0.d = 7'b0000001;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_cstopq48_nf_reg.d0_0 value=11 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_cstopq48_nf_reg.d0_0.d = 2'b11;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_efcnt_reg.d0_0 value=100100000000001 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_efcnt_reg.d0_0.d = 15'b100100000000001;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_efctl_reg.d0_0 value=111000 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_efctl_reg.d0_0.d = 6'b111000;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_enstat_reg.d0_0 value=1111111101111 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_enstat_reg.d0_0.d = 13'b1111111101111;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_flushclkstop_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_flushclkstop_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_foffcnt_nf_reg.d0_0 value=1101011 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_foffcnt_nf_reg.d0_0.d = 7'b1101011;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_fsreq_reg.d0_0 value=1 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_fsreq_reg.d0_0.d = 1'b1;

// instance=tb_top.cpu.tcu.sigmux_ctl.tcusig_rstsm_nf_reg.d0_0 value=01 out=q in=d model=dff 
force tb_top.cpu.tcu.sigmux_ctl.tcusig_rstsm_nf_reg.d0_0.d = 2'b01;


// 6260 forces installed

// Advance. Bench should be before posedge when this runs!
// For FC, lets try holding the forces for one cycle of the slowest
// clock and then release the forces.
// the release should be 38 clocks before the NCU unparks a thread.
@(posedge tb_top.SYSCLK);
@(negedge tb_top.SYSCLK);
#5; // exact time not critical

release tb_top.cpu.ccx.clk_ccx.xcluster_header_left.alatch.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_left.blatch_divr.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_left.ccu_div_ph_flop.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_left.clk_stopper.blatch.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_left.observe_flops.obs_ff2.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.alatch.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.blatch_divr.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.ccu_div_ph_flop.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.clk_stopper.blatch.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.ccx.clk_ccx.xcluster_header_right.observe_flops.obs_ff2.d;
release tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.cpx.bfd_io.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl0.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl1.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl2.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl3.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl4.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl5.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl6.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbl7.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr0.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr1.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr2.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr3.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr4.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr5.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr6.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.cpx.cpx_arbr7.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd0.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd0.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd0.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd0.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd1.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd1.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd1.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd1.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd2.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd2.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd2.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd2.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd3.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd3.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd3.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd3.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd4.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd4.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd4.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd4.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd5.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd5.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd5.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd5.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd6.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd6.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd6.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd6.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd7.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd7.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd7.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd7.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_0.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_1.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_2.d0_0.d;
release tb_top.cpu.ccx.pcx.bfd_io.i_dff_data_3.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl0.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl1.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl2.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl3.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl4.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl5.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl6.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl7.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbl8.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr0.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr1.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr2.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr3.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr4.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr5.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr6.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr7.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.dff_inreg_select.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q0.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q1.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q2.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q3.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q4.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q5.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q6.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q7.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.arc.q8.dff_qfullbar_a.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.ard.i_dff_qual_atomic_d1.d0_0.d;
release tb_top.cpu.ccx.pcx.pcx_arbr8.ard.i_dff_req_a.d0_0.d;
release tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.alatch.d;
release tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.blatch_divr.d;
release tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.dbg0.db0_clk_header_cmp_clk.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.dbg0.db0_clk_header_iol2clk.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.dbg0.rtc.ff_io_sync_en.d0_0.d;
release tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.alatch.d;
release tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.blatch_divr.d;
release tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.dbg1.db1_clk_header_cmp_clk.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.dbg1.db1_clk_header_iol2clk.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.dbg1.dbg1_dbgprt.ff_cmp_io_sync_en.d0_0.d;
release tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_0.d0_0.d;
release tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_1.d0_0.d;
release tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_data_2.d0_0.d;
release tb_top.cpu.dbg1.dbg1_dbgprt.ff_train_seq_gen.d0_0.d;
release tb_top.cpu.efu.efu_ioclk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.efu.efu_ioclk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.efu.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.efu.niu_interface.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.efu.niu_interface.ff_mcu_fclrz.d0_0.d;
release tb_top.cpu.efu.niu_interface.ff_niu_fclrz.d0_0.d;
release tb_top.cpu.efu.niu_interface.ff_psr_fclrz.d0_0.d;
release tb_top.cpu.efu.u_efa_stdc.enable_efa_por_reg.d0_0.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b0.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b0.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b0.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b0.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b0.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b0.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b0.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b0.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b0.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b0.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b0.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b0.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b0.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b0.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b0.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b0.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b0.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b0.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b0.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b1.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b1.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b1.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b1.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b1.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b1.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b1.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b1.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b1.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b1.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b1.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b1.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b1.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b1.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b1.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b1.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b1.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b1.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b1.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b2.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b2.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b2.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b2.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b2.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b2.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b2.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b2.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b2.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b2.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b2.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b2.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b2.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b2.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b2.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b2.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b2.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b2.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b2.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b3.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b3.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b3.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b3.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b3.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b3.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b3.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b3.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b3.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b3.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b3.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b3.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b3.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b3.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b3.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b3.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b3.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b3.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b3.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b4.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b4.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b4.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b4.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b4.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b4.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b4.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b4.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b4.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b4.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b4.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b4.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b4.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b4.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b4.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b4.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b4.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b4.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b4.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b5.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b5.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b5.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b5.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b5.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b5.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b5.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b5.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b5.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b5.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b5.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b5.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b5.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b5.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b5.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b5.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b5.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b5.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b5.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b6.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b6.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b6.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b6.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b6.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b6.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b6.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b6.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b6.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b6.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b6.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b6.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b6.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b6.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b6.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b6.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b6.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b6.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b6.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.alatch.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2b7.clock_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2b7.evict.ff_evict_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b7.evict.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b7.evict.ff_mux_select0_2b.d0_0.d;
release tb_top.cpu.l2b7.evict.ff_mux_select1_2a.d0_0.d;
release tb_top.cpu.l2b7.evict.ff_mux_select2_1b.d0_0.d;
release tb_top.cpu.l2b7.evict.ff_mux_select3_1a.d0_0.d;
release tb_top.cpu.l2b7.evict.ff_rdma_control_regs_slice.d0_0.d;
release tb_top.cpu.l2b7.fb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.fb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.fb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.fb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.fbd.ff_fb_rw_fail.d0_0.d;
release tb_top.cpu.l2b7.fbd.ff_fillbf_control_reg_slice.d0_0.d;
release tb_top.cpu.l2b7.l2d_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2b7.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2b7.rdma_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.rdma_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.rdma_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.rdma_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.rdmard.ff_sel_l1_slice.d0_0.d;
release tb_top.cpu.l2b7.rdmard.ff_sel_l2_slice.d0_0.d;
release tb_top.cpu.l2b7.rdmard.ff_sel_r1_slice.d0_0.d;
release tb_top.cpu.l2b7.rdmard.ff_sel_r2_slice.d0_0.d;
release tb_top.cpu.l2b7.rdmard.ff_select_inputs.d0_0.d;
release tb_top.cpu.l2b7.wb_array1.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.wb_array2.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.wb_array3.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2b7.wb_array4.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d0.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d0.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d0.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d0.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d0.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d0.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d0.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d0.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d0.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d1.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d1.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d1.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d1.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d1.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d1.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d1.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d1.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d1.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d2.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d2.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d2.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d2.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d2.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d2.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d2.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d2.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d2.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d3.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d3.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d3.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d3.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d3.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d3.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d3.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d3.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d3.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d4.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d4.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d4.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d4.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d4.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d4.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d4.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d4.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d4.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d5.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d5.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d5.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d5.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d5.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d5.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d5.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d5.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d5.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d6.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d6.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d6.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d6.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d6.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d6.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d6.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d6.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d6.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c4.d0_0.d;
release tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_00.d0_0.d;
release tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_01.d0_0.d;
release tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_20.d0_0.d;
release tb_top.cpu.l2d7.ctr.ff_cache_cache_rd_wr_c5_21.d0_0.d;
release tb_top.cpu.l2d7.l2d_clk_header.alatch.d;
release tb_top.cpu.l2d7.l2d_clk_header.blatch_divr.d;
release tb_top.cpu.l2d7.l2d_clk_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2d7.l2d_clk_header.clk_stopper.blatch.d;
release tb_top.cpu.l2d7.l2d_clk_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2d7.perif_io.ff_fill_clk_en_ov_stg.d0_0.d;
release tb_top.cpu.l2d7.perif_io.ff_l2t_l2d_rd_wr_c3.d0_0.d;
release tb_top.cpu.l2d7.perif_io.ff_pwrsav_ov_stg.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t0.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t0.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t0.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t0.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t0.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t0.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t0.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t0.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t0.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t0.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t0.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t0.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t0.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t0.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t0.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t0.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t0.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t0.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t0.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t0.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t0.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t0.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t0.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t0.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t0.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t0.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t0.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t0.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t0.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t0.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t0.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t0.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t0.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t0.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t0.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t0.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t0.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t0.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t0.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t0.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t0.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t0.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t0.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t0.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t0.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t0.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t0.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t0.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t0.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t0.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t0.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t0.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t0.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t0.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t0.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t0.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t0.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t0.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t0.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t0.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t0.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t0.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t0.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t0.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t0.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t0.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t0.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t0.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t0.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t0.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t0.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t0.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t0.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t0.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t0.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t0.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t0.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t0.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t0.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t0.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t0.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t0.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t0.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t0.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t0.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t0.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t0.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t0.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t0.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t0.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t0.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t0.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t0.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t0.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t0.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t0.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t0.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t0.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t1.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t1.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t1.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t1.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t1.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t1.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t1.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t1.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t1.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t1.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t1.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t1.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t1.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t1.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t1.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t1.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t1.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t1.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t1.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t1.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t1.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t1.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t1.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t1.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t1.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t1.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t1.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t1.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t1.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t1.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t1.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t1.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t1.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t1.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t1.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t1.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t1.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t1.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t1.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t1.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t1.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t1.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t1.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t1.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t1.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t1.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t1.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t1.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t1.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t1.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t1.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t1.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t1.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t1.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t1.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t1.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t1.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t1.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t1.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t1.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t1.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t1.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t1.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t1.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t1.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t1.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t1.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t1.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t1.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t1.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t1.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t1.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t1.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t1.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t1.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t1.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t1.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t1.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t1.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t1.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t1.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t1.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t1.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t1.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t1.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t1.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t1.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t1.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t1.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t1.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t1.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t1.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t1.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t1.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t1.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t1.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t1.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t1.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t2.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t2.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t2.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t2.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t2.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t2.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t2.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t2.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t2.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t2.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t2.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t2.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t2.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t2.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t2.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t2.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t2.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t2.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t2.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t2.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t2.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t2.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t2.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t2.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t2.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t2.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t2.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t2.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t2.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t2.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t2.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t2.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t2.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t2.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t2.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t2.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t2.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t2.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t2.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t2.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t2.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t2.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t2.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t2.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t2.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t2.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t2.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t2.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t2.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t2.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t2.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t2.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t2.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t2.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t2.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t2.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t2.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t2.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t2.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t2.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t2.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t2.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t2.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t2.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t2.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t2.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t2.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t2.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t2.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t2.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t2.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t2.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t2.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t2.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t2.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t2.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t2.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t2.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t2.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t2.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t2.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t2.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t2.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t2.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t2.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t2.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t2.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t2.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t2.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t2.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t2.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t2.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t2.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t2.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t2.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t2.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t2.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t2.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t3.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t3.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t3.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t3.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t3.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t3.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t3.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t3.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t3.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t3.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t3.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t3.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t3.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t3.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t3.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t3.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t3.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t3.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t3.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t3.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t3.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t3.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t3.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t3.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t3.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t3.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t3.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t3.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t3.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t3.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t3.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t3.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t3.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t3.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t3.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t3.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t3.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t3.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t3.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t3.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t3.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t3.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t3.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t3.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t3.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t3.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t3.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t3.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t3.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t3.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t3.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t3.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t3.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t3.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t3.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t3.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t3.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t3.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t3.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t3.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t3.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t3.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t3.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t3.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t3.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t3.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t3.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t3.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t3.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t3.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t3.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t3.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t3.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t3.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t3.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t3.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t3.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t3.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t3.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t3.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t3.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t3.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t3.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t3.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t3.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t3.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t3.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t3.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t3.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t3.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t3.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t3.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t3.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t3.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t3.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t3.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t3.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t3.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t4.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t4.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t4.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t4.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t4.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t4.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t4.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t4.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t4.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t4.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t4.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t4.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t4.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t4.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t4.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t4.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t4.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t4.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t4.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t4.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t4.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t4.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t4.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t4.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t4.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t4.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t4.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t4.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t4.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t4.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t4.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t4.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t4.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t4.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t4.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t4.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t4.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t4.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t4.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t4.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t4.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t4.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t4.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t4.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t4.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t4.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t4.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t4.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t4.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t4.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t4.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t4.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t4.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t4.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t4.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t4.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t4.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t4.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t4.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t4.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t4.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t4.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t4.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t4.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t4.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t4.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t4.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t4.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t4.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t4.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t4.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t4.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t4.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t4.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t4.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t4.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t4.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t4.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t4.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t4.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t4.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t4.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t4.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t4.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t4.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t4.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t4.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t4.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t4.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t4.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t4.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t4.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t4.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t4.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t4.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t4.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t4.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t4.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t5.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t5.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t5.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t5.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t5.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t5.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t5.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t5.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t5.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t5.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t5.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t5.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t5.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t5.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t5.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t5.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t5.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t5.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t5.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t5.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t5.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t5.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t5.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t5.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t5.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t5.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t5.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t5.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t5.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t5.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t5.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t5.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t5.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t5.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t5.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t5.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t5.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t5.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t5.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t5.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t5.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t5.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t5.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t5.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t5.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t5.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t5.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t5.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t5.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t5.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t5.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t5.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t5.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t5.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t5.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t5.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t5.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t5.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t5.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t5.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t5.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t5.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t5.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t5.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t5.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t5.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t5.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t5.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t5.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t5.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t5.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t5.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t5.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t5.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t5.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t5.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t5.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t5.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t5.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t5.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t5.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t5.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t5.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t5.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t5.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t5.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t5.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t5.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t5.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t5.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t5.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t5.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t5.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t5.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t5.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t5.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t5.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t5.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t6.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t6.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t6.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t6.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t6.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t6.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t6.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t6.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t6.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t6.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t6.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t6.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t6.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t6.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t6.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t6.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t6.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t6.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t6.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t6.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t6.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t6.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t6.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t6.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t6.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t6.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t6.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t6.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t6.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t6.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t6.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t6.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t6.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t6.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t6.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t6.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t6.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t6.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t6.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t6.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t6.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t6.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t6.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t6.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t6.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t6.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t6.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t6.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t6.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t6.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t6.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t6.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t6.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t6.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t6.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t6.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t6.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t6.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t6.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t6.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t6.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t6.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t6.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t6.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t6.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t6.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t6.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t6.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t6.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t6.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t6.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t6.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t6.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t6.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t6.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t6.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t6.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t6.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t6.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t6.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t6.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t6.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t6.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t6.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t6.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t6.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t6.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t6.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t6.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t6.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t6.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t6.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t6.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t6.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t6.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t6.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t6.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t6.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_arb_decdp_cas1_inst_c3.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_data_ecc_active_c4_dup.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_decdp_camld_inst_c2.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_decdp_ld_inst_c2.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_dword_mask_c8.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_ic_hitqual_cam_en_c3.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_parerr_gate_c1.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_waysel_gate_c2.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_word_lower_cmp_c9.d0_0.d;
release tb_top.cpu.l2t7.arb.ff_word_upper_cmp_c9.d0_0.d;
release tb_top.cpu.l2t7.arb.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.arbadr.ff_mux3_bufsel_px2.d0_0.d;
release tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_1.d0_0.d;
release tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_2.d0_0.d;
release tb_top.cpu.l2t7.arbadr.ff_ncu_mux_sel_3.d0_0.d;
release tb_top.cpu.l2t7.arbadr.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t7.arbdat.ff_col_offset_sel_c2.d0_0.d;
release tb_top.cpu.l2t7.arbdat.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t7.arbdec.ff_inst_size_c8.d0_0.d;
release tb_top.cpu.l2t7.arbdec.ff_mbdata_mbist_reg.d0_0.d;
release tb_top.cpu.l2t7.csreg.ff_mux1_sel_c7.d0_0.d;
release tb_top.cpu.l2t7.dc_out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.dc_out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.dc_out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.dc_out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.dc_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.dc_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t7.dc_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t7.dc_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t7.dc_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.dc_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.dc_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t7.dc_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t7.dc_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t7.dc_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t7.decc.ff_fame_mbist_flops_0.d0_0.d;
release tb_top.cpu.l2t7.deccck.ff_deccck_muxsel_diag_out_c7.d0_0.d;
release tb_top.cpu.l2t7.dirrep.ff_dir_vld_dcd_c4_l.d0_0.d;
release tb_top.cpu.l2t7.dirrep.ff_inval_mask_dcd_c4.d0_0.d;
release tb_top.cpu.l2t7.dirrep.ff_inval_mask_icd_c4.d0_0.d;
release tb_top.cpu.l2t7.dirvec.ff_ncu_signals.d0_0.d;
release tb_top.cpu.l2t7.dirvec.ff_staged_part_bank.d0_0.d;
release tb_top.cpu.l2t7.dirvec.ff_sync_en.d0_0.d;
release tb_top.cpu.l2t7.dmologic.ff_dmo_data_1.d0_0.d;
release tb_top.cpu.l2t7.evctag.ff_shifted_index.d0_0.d;
release tb_top.cpu.l2t7.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t7.fbtag.xx62.d0_0.d;
release tb_top.cpu.l2t7.filbuf.ff_fb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t7.filbuf.ff_fill_entry_num_c2.d0_0.d;
release tb_top.cpu.l2t7.filbuf.ff_fill_entry_num_c3.d0_0.d;
release tb_top.cpu.l2t7.filbuf.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t7.filbuf.ff_l2_rd_state.d0_0.d;
release tb_top.cpu.l2t7.filbuf.ff_l2_rd_state_quad0.d0_0.d;
release tb_top.cpu.l2t7.filbuf.ff_l2_rd_state_quad1.d0_0.d;
release tb_top.cpu.l2t7.filbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.ic_row0.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.ic_row0.wr_data0_so_15.d;
release tb_top.cpu.l2t7.ic_row0.wr_data1_so_15.d;
release tb_top.cpu.l2t7.ic_row0.wr_data2_so_15.d;
release tb_top.cpu.l2t7.ic_row0.wr_data3_so_15.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask0_so_7.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask1_so_7.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask2_so_7.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_0.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_1.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_2.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_3.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_4.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_5.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_6.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.ic_row2.inv_mask3_so_7.d;
release tb_top.cpu.l2t7.ic_row2.wr_data0_so_15.d;
release tb_top.cpu.l2t7.ic_row2.wr_data1_so_15.d;
release tb_top.cpu.l2t7.ic_row2.wr_data2_so_15.d;
release tb_top.cpu.l2t7.ic_row2.wr_data3_so_15.d;
release tb_top.cpu.l2t7.iqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t7.iqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.iqu.ff_array_wr_ptr_plus1.d0_0.d;
release tb_top.cpu.l2t7.iqu.ff_iqu_sel_pcx.d0_0.d;
release tb_top.cpu.l2t7.iqu.ff_que_cnt_0.d0_0.d;
release tb_top.cpu.l2t7.iqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.ique.ff_pcx_l2t_data_c1_2.d0_0.d;
release tb_top.cpu.l2t7.l2drpt.ff_all_signals.d0_0.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.alatch.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.blatch_divr.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.l2t7.l2t_clk_header.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.l2t7.l2tag_sram_hdr.efuse_l2d_header.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.l2t7.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t7.mb2_control.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t7.mbdata.ff_wdata_1.d0_0.d;
release tb_top.cpu.l2t7.mbist.input_signals_reg.d0_0.d;
release tb_top.cpu.l2t7.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t7.mbtag.xx84.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_fbsel_def_vld_d1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_idx_c1c2comp_c1_d1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad0.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad2.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad3.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad4.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad5.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad6.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_l2_state_quad7.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mb_hit_off_c1_d1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mb_write_ptr_c3.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c4.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c5.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c52.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c6.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c7.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mbf_dep_c8.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_pick_2_l.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad0.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad2.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad3.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad4.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad5.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad6.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_mcu_state_quad7.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_misbuf_c1c2_match_c1_d1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_misbuf_c1c2_match_c1_d1_1.d0_0.d;
release tb_top.cpu.l2t7.misbuf.ff_set_dep_c2_ldifetch_miss_c2.d0_0.d;
release tb_top.cpu.l2t7.misbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.oqarray.ff_byte_wen.d0_0.d;
release tb_top.cpu.l2t7.oqarray.ff_wdata_72.d0_0.d;
release tb_top.cpu.l2t7.oqarray.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_allow_req_c7.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_dec_cpu_c52.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_dec_cpu_c6.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_dec_cpu_c7.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_dec_cpuid_c6.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_diag_def_sel_c8.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_mux_vec_sel_c52.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_mux_vec_sel_c6.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_oq_cnt_minus1_d1.d0_0.d;
release tb_top.cpu.l2t7.oqu.ff_oq_cnt_plus1_d1.d0_0.d;
release tb_top.cpu.l2t7.oqu.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.oque.ff_data_rtn_d1_1.d0_0.d;
release tb_top.cpu.l2t7.oque.ff_mbist_flop.d0_0.d;
release tb_top.cpu.l2t7.oque.ff_tmp_cpx_data_ca_1.d0_0.d;
release tb_top.cpu.l2t7.out_col0.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.out_col1.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.out_col2.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.out_col3.ff_lookup_cmp_data.d0_0.d;
release tb_top.cpu.l2t7.rdmat.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t7.rdmat.ff_rdma_wr_ptr_s2.d0_0.d;
release tb_top.cpu.l2t7.rdmat.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t7.rdmatag.xx62.d0_0.d;
release tb_top.cpu.l2t7.snp.ff_snp_rdmatag_wr_en_s2_4muxsel_d1.d0_0.d;
release tb_top.cpu.l2t7.snp.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.snpd.ff_snp_rd_ptr_d1_5_MERGED.d0_0.d;
release tb_top.cpu.l2t7.subarray_0.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.subarray_1.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.subarray_10.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.subarray_11.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.subarray_2.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.subarray_3.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.subarray_8.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.subarray_9.ff_word_wen.d0_0.d;
release tb_top.cpu.l2t7.tag.ff_clk_en_ov.d0_0.d;
release tb_top.cpu.l2t7.tag.ff_ff_wr_en_ov.d0_0.d;
release tb_top.cpu.l2t7.tag.quad0.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad0.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tag.quad0.bank0.reg_wr_way_b.d0_0.d;
release tb_top.cpu.l2t7.tag.quad0.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad0.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tag.quad1.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad1.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tag.quad1.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad1.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tag.quad2.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad2.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tag.quad2.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad2.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tag.quad3.bank0.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad3.bank0.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tag.quad3.bank1.reg_way_hit_a0.d0_0.d;
release tb_top.cpu.l2t7.tag.quad3.bank1.reg_way_hit_a1.d0_0.d;
release tb_top.cpu.l2t7.tagctl.ff_alt_tag_miss_unqual_c3.d0_0.d;
release tb_top.cpu.l2t7.tagctl.ff_l2_bypass_mode_on.d0_0.d;
release tb_top.cpu.l2t7.tagctl.ff_ld_inst_c3.d0_0.d;
release tb_top.cpu.l2t7.tagctl.ff_prev_wen_c1.d0_0.d;
release tb_top.cpu.l2t7.tagctl.ff_scrub_wr_disable_c9.d0_0.d;
release tb_top.cpu.l2t7.tagctl.ff_tag_l2b_fbd_stdatasel_c3.d0_0.d;
release tb_top.cpu.l2t7.tagctl.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.tagd.ff_ecc_staging5_8.d0_0.d;
release tb_top.cpu.l2t7.tagd.ff_piped_vuad0.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_dir_quad_way_c3.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_quad_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_state.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_state_quad0.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_state_quad1.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_state_quad2.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_state_quad3.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_way_c3.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_lru_way_c3_1.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_tag_quad0_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_tag_quad1_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_tag_quad2_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_tag_quad3_muxsel_c2.d0_0.d;
release tb_top.cpu.l2t7.tagdp.ff_use_dec_sel_c3.d0_0.d;
release tb_top.cpu.l2t7.tagdp.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.usaloc.ff_used_alloc_c3.d0_0.d;
release tb_top.cpu.l2t7.usaloc.ff_used_and_alloc_rd_c2.d0_0.d;
release tb_top.cpu.l2t7.vlddir.ff_valid_dirty_rd_c2.d0_0.d;
release tb_top.cpu.l2t7.vuad.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t7.vuad.ff_vuaddp_vuad_sel_c2.d0_0.d;
release tb_top.cpu.l2t7.vuadpm.ff_mbist_write_data.d0_0.d;
release tb_top.cpu.l2t7.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t7.wbtag.xx62.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_arb_wbuf_hit_off_c2.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_l2_bypass_mode_on_d1.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_quad0_state.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_quad1_state.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_quad2_state.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_quad_state.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_state.d0_0.d;
release tb_top.cpu.l2t7.wbuf.ff_wbtag_write_wl_c5.d0_0.d;
release tb_top.cpu.l2t7.wbuf.reset_flop.d0_0.d;
release tb_top.cpu.l2t7.wbufrpt.ff_l2t_l2b_evict_en_r0.d0_0.d;
release tb_top.cpu.mcu0.clkgen_cmp.xcluster_header.alatch.d;
release tb_top.cpu.mcu0.clkgen_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu0.clkgen_dr.xcluster_header.alatch.d;
release tb_top.cpu.mcu0.clkgen_dr.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu0.clkgen_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu0.drif.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu0.drif.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu0.drif.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu0.drif.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu0.drif.ff_dal_reg.d0_0.d;
release tb_top.cpu.mcu0.drif.ff_err_fifo_empty_d1.d0_0.d;
release tb_top.cpu.mcu0.drif.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu0.drif.ff_ral_reg.d0_0.d;
release tb_top.cpu.mcu0.drif.ff_sync_frame_req_l.d0_0.d;
release tb_top.cpu.mcu0.drif.ff_time_cntr.d0_0.d;
release tb_top.cpu.mcu0.drif.reqq.woq.ff_io_wdata_sel.d0_0.d;
release tb_top.cpu.mcu0.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_chnl_latency_cntr.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_config_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_crc_sel0.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_crc_sel1.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_elect_idle_detect.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_l0s_stall.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_polling_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_tclktrain_min_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_tclktrain_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_tdisable_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_testing_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_ts_match0.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_ts_match0_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_ts_match1.d0_0.d;
release tb_top.cpu.mcu0.fbdic.ff_ts_match1_cnt.d0_0.d;
release tb_top.cpu.mcu0.fbdic.spare20_flop.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll0.xx0.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll0.xx1.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll1.xx0.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll1.xx1.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll2.xx0.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll2.xx1.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll3.xx0.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll3.xx1.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll4.xx0.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll4.xx1.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll5.xx0.d;
release tb_top.cpu.mcu0.fbdic.sync_stspll5.xx1.d;
release tb_top.cpu.mcu0.fdoklu.ff_idle_lfsr.d0_0.d;
release tb_top.cpu.mcu0.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d;
release tb_top.cpu.mcu0.fdout.spare0_flop.d;
release tb_top.cpu.mcu0.l2if0.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu0.l2if0.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu0.l2if0.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu0.l2if0.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu0.l2if0.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu0.l2if0.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu0.l2if0.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu0.l2if1.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu0.l2if1.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu0.l2if1.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu0.l2if1.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu0.l2if1.ff_addr.d0_0.d;
release tb_top.cpu.mcu0.l2if1.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu0.l2if1.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu0.l2if1.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu0.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu0.mbist.data_pipe_reg1.d0_0.d;
release tb_top.cpu.mcu0.mbist.data_pipe_reg2.d0_0.d;
release tb_top.cpu.mcu0.mbist.data_pipe_reg3.d0_0.d;
release tb_top.cpu.mcu0.mbist.data_pipe_reg4.d0_0.d;
release tb_top.cpu.mcu0.mbist.wdata_reg.d0_0.d;
release tb_top.cpu.mcu0.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d;
release tb_top.cpu.mcu0.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d;
release tb_top.cpu.mcu0.rdata.ff_io_sync_pulses.d0_0.d;
release tb_top.cpu.mcu0.rdata.ff_mbist_data.d0_0.d;
release tb_top.cpu.mcu0.rdata.ff_mcu_sync_pulse_delays.d0_0.d;
release tb_top.cpu.mcu0.rdata.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu0.rdata.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu0.ucb.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu0.wrdp.u_io_ecc_15_0.d0_0.d;
release tb_top.cpu.mcu1.clkgen_cmp.xcluster_header.alatch.d;
release tb_top.cpu.mcu1.clkgen_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu1.clkgen_dr.xcluster_header.alatch.d;
release tb_top.cpu.mcu1.clkgen_dr.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu1.clkgen_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu1.drif.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu1.drif.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu1.drif.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu1.drif.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu1.drif.ff_dal_reg.d0_0.d;
release tb_top.cpu.mcu1.drif.ff_err_fifo_empty_d1.d0_0.d;
release tb_top.cpu.mcu1.drif.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu1.drif.ff_ral_reg.d0_0.d;
release tb_top.cpu.mcu1.drif.ff_sync_frame_req_l.d0_0.d;
release tb_top.cpu.mcu1.drif.ff_time_cntr.d0_0.d;
release tb_top.cpu.mcu1.drif.reqq.woq.ff_io_wdata_sel.d0_0.d;
release tb_top.cpu.mcu1.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_chnl_latency_cntr.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_config_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_crc_sel0.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_crc_sel1.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_elect_idle_detect.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_l0s_stall.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_polling_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_tclktrain_min_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_tclktrain_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_tdisable_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_testing_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_ts_match0.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_ts_match0_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_ts_match1.d0_0.d;
release tb_top.cpu.mcu1.fbdic.ff_ts_match1_cnt.d0_0.d;
release tb_top.cpu.mcu1.fbdic.spare20_flop.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll0.xx0.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll0.xx1.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll1.xx0.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll1.xx1.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll2.xx0.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll2.xx1.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll3.xx0.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll3.xx1.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll4.xx0.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll4.xx1.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll5.xx0.d;
release tb_top.cpu.mcu1.fbdic.sync_stspll5.xx1.d;
release tb_top.cpu.mcu1.fdoklu.ff_idle_lfsr.d0_0.d;
release tb_top.cpu.mcu1.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d;
release tb_top.cpu.mcu1.fdout.spare0_flop.d;
release tb_top.cpu.mcu1.l2if0.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu1.l2if0.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu1.l2if0.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu1.l2if0.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu1.l2if0.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu1.l2if0.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu1.l2if0.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu1.l2if1.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu1.l2if1.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu1.l2if1.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu1.l2if1.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu1.l2if1.ff_addr.d0_0.d;
release tb_top.cpu.mcu1.l2if1.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu1.l2if1.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu1.l2if1.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu1.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu1.mbist.data_pipe_reg1.d0_0.d;
release tb_top.cpu.mcu1.mbist.data_pipe_reg2.d0_0.d;
release tb_top.cpu.mcu1.mbist.data_pipe_reg3.d0_0.d;
release tb_top.cpu.mcu1.mbist.data_pipe_reg4.d0_0.d;
release tb_top.cpu.mcu1.mbist.wdata_reg.d0_0.d;
release tb_top.cpu.mcu1.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d;
release tb_top.cpu.mcu1.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d;
release tb_top.cpu.mcu1.rdata.ff_io_sync_pulses.d0_0.d;
release tb_top.cpu.mcu1.rdata.ff_mbist_data.d0_0.d;
release tb_top.cpu.mcu1.rdata.ff_mcu_sync_pulse_delays.d0_0.d;
release tb_top.cpu.mcu1.rdata.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu1.rdata.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu1.ucb.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu1.wrdp.u_io_ecc_15_0.d0_0.d;
release tb_top.cpu.mcu2.clkgen_cmp.xcluster_header.alatch.d;
release tb_top.cpu.mcu2.clkgen_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu2.clkgen_dr.xcluster_header.alatch.d;
release tb_top.cpu.mcu2.clkgen_dr.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu2.clkgen_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu2.drif.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu2.drif.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu2.drif.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu2.drif.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu2.drif.ff_dal_reg.d0_0.d;
release tb_top.cpu.mcu2.drif.ff_err_fifo_empty_d1.d0_0.d;
release tb_top.cpu.mcu2.drif.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu2.drif.ff_ral_reg.d0_0.d;
release tb_top.cpu.mcu2.drif.ff_sync_frame_req_l.d0_0.d;
release tb_top.cpu.mcu2.drif.ff_time_cntr.d0_0.d;
release tb_top.cpu.mcu2.drif.reqq.woq.ff_io_wdata_sel.d0_0.d;
release tb_top.cpu.mcu2.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_chnl_latency_cntr.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_config_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_crc_sel0.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_crc_sel1.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_elect_idle_detect.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_l0s_stall.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_polling_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_tclktrain_min_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_tclktrain_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_tdisable_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_testing_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_ts_match0.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_ts_match0_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_ts_match1.d0_0.d;
release tb_top.cpu.mcu2.fbdic.ff_ts_match1_cnt.d0_0.d;
release tb_top.cpu.mcu2.fbdic.spare20_flop.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll0.xx0.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll0.xx1.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll1.xx0.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll1.xx1.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll2.xx0.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll2.xx1.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll3.xx0.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll3.xx1.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll4.xx0.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll4.xx1.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll5.xx0.d;
release tb_top.cpu.mcu2.fbdic.sync_stspll5.xx1.d;
release tb_top.cpu.mcu2.fdoklu.ff_idle_lfsr.d0_0.d;
release tb_top.cpu.mcu2.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d;
release tb_top.cpu.mcu2.fdout.spare0_flop.d;
release tb_top.cpu.mcu2.l2if0.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu2.l2if0.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu2.l2if0.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu2.l2if0.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu2.l2if0.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu2.l2if0.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu2.l2if0.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu2.l2if1.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu2.l2if1.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu2.l2if1.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu2.l2if1.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu2.l2if1.ff_addr.d0_0.d;
release tb_top.cpu.mcu2.l2if1.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu2.l2if1.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu2.l2if1.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu2.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu2.mbist.data_pipe_reg1.d0_0.d;
release tb_top.cpu.mcu2.mbist.data_pipe_reg2.d0_0.d;
release tb_top.cpu.mcu2.mbist.data_pipe_reg3.d0_0.d;
release tb_top.cpu.mcu2.mbist.data_pipe_reg4.d0_0.d;
release tb_top.cpu.mcu2.mbist.wdata_reg.d0_0.d;
release tb_top.cpu.mcu2.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d;
release tb_top.cpu.mcu2.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d;
release tb_top.cpu.mcu2.rdata.ff_io_sync_pulses.d0_0.d;
release tb_top.cpu.mcu2.rdata.ff_mbist_data.d0_0.d;
release tb_top.cpu.mcu2.rdata.ff_mcu_sync_pulse_delays.d0_0.d;
release tb_top.cpu.mcu2.rdata.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu2.rdata.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu2.ucb.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu2.wrdp.u_io_ecc_15_0.d0_0.d;
release tb_top.cpu.mcu3.clkgen_cmp.xcluster_header.alatch.d;
release tb_top.cpu.mcu3.clkgen_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu3.clkgen_dr.xcluster_header.alatch.d;
release tb_top.cpu.mcu3.clkgen_dr.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu3.clkgen_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mcu3.drif.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu3.drif.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu3.drif.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu3.drif.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu3.drif.ff_dal_reg.d0_0.d;
release tb_top.cpu.mcu3.drif.ff_err_fifo_empty_d1.d0_0.d;
release tb_top.cpu.mcu3.drif.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu3.drif.ff_ral_reg.d0_0.d;
release tb_top.cpu.mcu3.drif.ff_sync_frame_req_l.d0_0.d;
release tb_top.cpu.mcu3.drif.ff_time_cntr.d0_0.d;
release tb_top.cpu.mcu3.drif.reqq.woq.ff_io_wdata_sel.d0_0.d;
release tb_top.cpu.mcu3.fbdic.fbdtm.ff_idle_lfsr_reset.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_chnl_latency_cntr.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_config_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_crc_sel0.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_crc_sel1.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_elect_idle_detect.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_l0s_stall.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_polling_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_tclktrain_min_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_tclktrain_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_tdisable_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_testing_timeout_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_ts_match0.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_ts_match0_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_ts_match1.d0_0.d;
release tb_top.cpu.mcu3.fbdic.ff_ts_match1_cnt.d0_0.d;
release tb_top.cpu.mcu3.fbdic.spare20_flop.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll0.xx0.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll0.xx1.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll1.xx0.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll1.xx1.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll2.xx0.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll2.xx1.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll3.xx0.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll3.xx1.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll4.xx0.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll4.xx1.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll5.xx0.d;
release tb_top.cpu.mcu3.fbdic.sync_stspll5.xx1.d;
release tb_top.cpu.mcu3.fdoklu.ff_idle_lfsr.d0_0.d;
release tb_top.cpu.mcu3.fdoklu.ff_link_cnt_eq_0_d1.d0_0.d;
release tb_top.cpu.mcu3.fdout.spare0_flop.d;
release tb_top.cpu.mcu3.l2if0.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu3.l2if0.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu3.l2if0.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu3.l2if0.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu3.l2if0.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu3.l2if0.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu3.l2if0.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu3.l2if1.adrgen.ff_error_mask.d0_0.d;
release tb_top.cpu.mcu3.l2if1.adrgen.ff_mem_type.d0_0.d;
release tb_top.cpu.mcu3.l2if1.adrgen.ff_num_dimms.d0_0.d;
release tb_top.cpu.mcu3.l2if1.adrgen.ff_rank_mask.d0_0.d;
release tb_top.cpu.mcu3.l2if1.ff_addr.d0_0.d;
release tb_top.cpu.mcu3.l2if1.ff_addr_mode.d0_0.d;
release tb_top.cpu.mcu3.l2if1.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu3.l2if1.ff_partial_mode.d0_0.d;
release tb_top.cpu.mcu3.l2rdmx.u_l2ecc_mbist_wdata.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw0.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf0.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf1.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf10.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf11.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf12.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf13.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf2.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf3.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf4.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf5.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf6.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf7.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf8.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.lndskw1.algnbf9.ff_rptr_wptr.d0_0.d;
release tb_top.cpu.mcu3.mbist.data_pipe_reg1.d0_0.d;
release tb_top.cpu.mcu3.mbist.data_pipe_reg2.d0_0.d;
release tb_top.cpu.mcu3.mbist.data_pipe_reg3.d0_0.d;
release tb_top.cpu.mcu3.mbist.data_pipe_reg4.d0_0.d;
release tb_top.cpu.mcu3.mbist.wdata_reg.d0_0.d;
release tb_top.cpu.mcu3.rdata.ff_ddr_cmp_sync_en_d12.d0_0.d;
release tb_top.cpu.mcu3.rdata.ff_ddr_cmp_sync_en_d23.d0_0.d;
release tb_top.cpu.mcu3.rdata.ff_io_sync_pulses.d0_0.d;
release tb_top.cpu.mcu3.rdata.ff_mbist_data.d0_0.d;
release tb_top.cpu.mcu3.rdata.ff_mcu_sync_pulse_delays.d0_0.d;
release tb_top.cpu.mcu3.rdata.ff_mcu_sync_pulses.d0_0.d;
release tb_top.cpu.mcu3.rdata.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu3.ucb.ff_partial_bank_mode.d0_0.d;
release tb_top.cpu.mcu3.wrdp.u_io_ecc_15_0.d0_0.d;
release tb_top.cpu.mio.cell_10.ff_in.d;
release tb_top.cpu.mio.cell_103.ff_in.d;
release tb_top.cpu.mio.cell_104.ff_in.d;
release tb_top.cpu.mio.cell_105.ff_in.d;
release tb_top.cpu.mio.cell_106.ff_in.d;
release tb_top.cpu.mio.cell_107.ff_in.d;
release tb_top.cpu.mio.cell_108.ff_in.d;
release tb_top.cpu.mio.cell_110.ff_in.d;
release tb_top.cpu.mio.cell_12.ff_in.d;
release tb_top.cpu.mio.cell_129.ff_in.d;
release tb_top.cpu.mio.cell_13.ff_in.d;
release tb_top.cpu.mio.cell_130.ff_in.d;
release tb_top.cpu.mio.cell_131.ff_in.d;
release tb_top.cpu.mio.cell_132.ff_in.d;
release tb_top.cpu.mio.cell_133.ff_in.d;
release tb_top.cpu.mio.cell_134.ff_in.d;
release tb_top.cpu.mio.cell_135.ff_in.d;
release tb_top.cpu.mio.cell_136.ff_in.d;
release tb_top.cpu.mio.cell_137.ff_in.d;
release tb_top.cpu.mio.cell_138.ff_in.d;
release tb_top.cpu.mio.cell_139.ff_in.d;
release tb_top.cpu.mio.cell_14.ff_in.d;
release tb_top.cpu.mio.cell_140.ff_in.d;
release tb_top.cpu.mio.cell_141.ff_in.d;
release tb_top.cpu.mio.cell_142.ff_in.d;
release tb_top.cpu.mio.cell_143.ff_in.d;
release tb_top.cpu.mio.cell_144.ff_in.d;
release tb_top.cpu.mio.cell_145.ff_in.d;
release tb_top.cpu.mio.cell_146.ff_in.d;
release tb_top.cpu.mio.cell_147.ff_in.d;
release tb_top.cpu.mio.cell_148.ff_in.d;
release tb_top.cpu.mio.cell_149.ff_in.d;
release tb_top.cpu.mio.cell_15.ff_oe.d;
release tb_top.cpu.mio.cell_15.ff_out.d;
release tb_top.cpu.mio.cell_150.ff_in.d;
release tb_top.cpu.mio.cell_151.ff_in.d;
release tb_top.cpu.mio.cell_152.ff_in.d;
release tb_top.cpu.mio.cell_153.ff_in.d;
release tb_top.cpu.mio.cell_154.ff_in.d;
release tb_top.cpu.mio.cell_155.ff_in.d;
release tb_top.cpu.mio.cell_156.ff_in.d;
release tb_top.cpu.mio.cell_157.ff_in.d;
release tb_top.cpu.mio.cell_158.ff_in.d;
release tb_top.cpu.mio.cell_159.ff_in.d;
release tb_top.cpu.mio.cell_160.ff_in.d;
release tb_top.cpu.mio.cell_161.ff_in.d;
release tb_top.cpu.mio.cell_162.ff_in.d;
release tb_top.cpu.mio.cell_163.ff_in.d;
release tb_top.cpu.mio.cell_164.ff_in.d;
release tb_top.cpu.mio.cell_165.ff_in.d;
release tb_top.cpu.mio.cell_17.ff_oe.d;
release tb_top.cpu.mio.cell_176.ff_in.d;
release tb_top.cpu.mio.cell_177.ff_in.d;
release tb_top.cpu.mio.cell_178.ff_in.d;
release tb_top.cpu.mio.cell_179.ff_in.d;
release tb_top.cpu.mio.cell_18.ff_oe.d;
release tb_top.cpu.mio.cell_180.ff_in.d;
release tb_top.cpu.mio.cell_181.ff_in.d;
release tb_top.cpu.mio.cell_182.ff_in.d;
release tb_top.cpu.mio.cell_184.ff_in.d;
release tb_top.cpu.mio.cell_186.ff_out.d;
release tb_top.cpu.mio.cell_187.ff_out.d;
release tb_top.cpu.mio.cell_189.ff_out.d;
release tb_top.cpu.mio.cell_193.ff_in.d;
release tb_top.cpu.mio.cell_2.ff_oe.d;
release tb_top.cpu.mio.cell_202.ff_oe.d;
release tb_top.cpu.mio.cell_209.ff_oe.d;
release tb_top.cpu.mio.cell_210.ff_oe.d;
release tb_top.cpu.mio.cell_211.ff_in.d;
release tb_top.cpu.mio.cell_211.ff_out.d;
release tb_top.cpu.mio.cell_23.ff_in.d;
release tb_top.cpu.mio.cell_24.ff_oe.d;
release tb_top.cpu.mio.cell_27.ff_in_mux_data.d0_0.d;
release tb_top.cpu.mio.cell_3.ff_oe.d;
release tb_top.cpu.mio.cell_3.ff_out.d;
release tb_top.cpu.mio.cell_4.ff_in.d;
release tb_top.cpu.mio.cell_5.ff_oe.d;
release tb_top.cpu.mio.cell_6.ff_oe.d;
release tb_top.cpu.mio.cell_7.ff_oe.d;
release tb_top.cpu.mio.cell_7.ff_out.d;
release tb_top.cpu.mio.cell_8.ff_in.d;
release tb_top.cpu.mio.cell_9.ff_oe.d;
release tb_top.cpu.mio.cell_9.ff_out.d;
release tb_top.cpu.mio.cell_98.ff_in.d;
release tb_top.cpu.mio.io2xsyncen_reg0.ff_0.d0_0.d;
release tb_top.cpu.mio.io2xsyncen_reg1.ff_0.d0_0.d;
release tb_top.cpu.mio.io2xsyncen_reg2.ff_0.d0_0.d;
release tb_top.cpu.mio.io2xsyncen_reg3.ff_0.d0_0.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.alatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.blatch_divr.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_0.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.alatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.blatch_divr.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_1.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.alatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.blatch_divr.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_2.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.alatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.blatch_divr.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mio.mio_clk_header_cmp_clk_3.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.mio.mio_clk_header_iol2clk.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.mio.muxsel.ff_1.d0_1.d;
release tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.alatch.d;
release tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.blatch_divr.d;
release tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.ncu.clkgen_ncu_cmp.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.ncu.clkgen_ncu_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.ncu.ncu_cpu_buf_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_cpu_buf_rf_cust.dff_dout.d0_0.d;
release tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_din_lo.d0_0.d;
release tb_top.cpu.ncu.ncu_dmubuf0_rf_cust.dff_dout.d0_0.d;
release tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_din_lo.d0_0.d;
release tb_top.cpu.ncu.ncu_dmubuf1_rf_cust.dff_dout.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.io_cmp_sync_en_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifc_ctl.cpu_mondo_addr_creg_mdata0_dec_d1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo2cpu_pkt_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_busy_dout_d2_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_busy_vec_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data0_din_d1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data0_din_d2_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data1_din_d1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_c2ifcd_ctl.ncu_c2ifd_ctl.mondo_data1_din_d2_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.intbuf_pa_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.iobuf_pa_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg1.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg2.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.data_pipe_reg3.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.mb0_wdata_reg.d0_0.d;
release tb_top.cpu.ncu.ncu_fcd_ctl.ncu_mb0_ctl.res_read_data_reg.d0_0.d;
release tb_top.cpu.ncu.ncu_intbuf_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_intbuf_rf_cust.dff_dout.d0_0.d;
release tb_top.cpu.ncu.ncu_intman_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_intman_rf_cust.dff_rd_en.d0_0.d;
release tb_top.cpu.ncu.ncu_intman_rf_cust.dff_rd_en.d0_0.d;
release tb_top.cpu.ncu.ncu_iobuf0_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_iobuf0_rf_cust.dff_dout.d0_0.d;
release tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_din_lo.d0_0.d;
release tb_top.cpu.ncu.ncu_iobuf1_rf_cust.dff_dout.d0_0.d;
release tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_rd_en.d0_0.d;
release tb_top.cpu.ncu.ncu_mondo0_rf_cust.dff_rd_en.d0_0.d;
release tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_din_hi.d0_0.d;
release tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_rd_en.d0_0.d;
release tb_top.cpu.ncu.ncu_mondo1_rf_cust.dff_rd_en.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ccu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ccu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dbg1_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dbg1_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmucsr_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmucsr_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.cr_id_rtn1_par_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.ncu_dmu_dpar_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.pad_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu0_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu0_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu1_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu1_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu2_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu2_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu3_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.mcu3_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_c2isd_ctl.cpubuf_pa_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.core_running_status0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.fusestat_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.l2pm_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.l2pm_preview_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_ctrl_ctl.por_upd_en_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg1.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg2.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg3.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.cmpsel_pipe_reg4.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg1.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg2.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.data_pipe_reg3.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.mb1_wdata_reg.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_mb1_ctl.res_read_data_reg.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.niu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.niu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.rcu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.rcu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ssi_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ssi_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.tcu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.tcu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ccu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ccu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dbg1_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dbg1_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dmucsr_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.dmucsr_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu0_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu0_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu1_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu1_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu2_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu2_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu3_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.mcu3_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ncu_i2csc_ctl.mondo_busy_d1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ncu_i2csc_ctl.mondo_busy_vec_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.niu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.niu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.rcu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.rcu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.ncu_dmu_mondo_id_par_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.sii_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ssi_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.ssi_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.tcu_ucb_buf.rdy0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_scd_ctl.ncu_i2cscd_ctl.tcu_ucb_buf.rdy1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.cntr_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.sck_cnt_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.sck_posedge_d3_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_async_ctu_jbi_ssiclk_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_async_jbi_io_ssi_sck.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dffrl_sck_cyc_cnt.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg3.p_out_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg4.p_out_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg5.p_out_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg6.p_out_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_mosi_shreg7.p_out_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.toreg_ld0_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.toreg_ld1_ff.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d1.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d2.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d3.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d4.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d5.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d6.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_ext_int_l_d7.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_io_jbi_ext_int_l_pre_sync.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_io_jbi_ext_int_l_sync.d0_0.d;
release tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssiuif_ctl.u_dff_timeout_reg.d0_0.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.alatch.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.blatch_divr.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.rst.clkgen_rst_cmp.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.rst.clkgen_rst_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.rst.clkgen_rst_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.rst.rst_cmp_ctl.ccu_rst_change_cmp0_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.ccu_rst_change_cmp_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.io_cmp_sync_en2_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.mio_rst_pb_rst_cmp_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.mio_rst_pb_rst_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_cmp_ctl_wmr_cmp_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_dmu_peu_por_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_dmu_peu_wmr_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_l2_por_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_l2_wmr_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_niu_mac_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_niu_wmr_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_rst_por_cmp_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_rst_por_io_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_rst_pwron_rst_l_io0_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_rst_wmr_cmp_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_rst_wmr_io_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.rst_tcu_pwron_rst_l_ff.d0_0.d;
release tb_top.cpu.rst.rst_cmp_ctl.tcu_rst_flush_stop_ack_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.ccu_count_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.ccu_rst_change_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.cluster_arst_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.lock_count_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.mio_rst_button_xir_sys_ff.xx0.d;
release tb_top.cpu.rst.rst_fsm_ctl.mio_rst_button_xir_sys_ff.xx1.d;
release tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys3_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys_ff.xx0.d;
release tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pb_rst_sys_ff.xx1.d;
release tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pwron_rst_sys_ff.xx0.d;
release tb_top.cpu.rst.rst_fsm_ctl.mio_rst_pwron_rst_sys_ff.xx1.d;
release tb_top.cpu.rst.rst_fsm_ctl.niu_count_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.prop_count_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_ccu_pll_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_ccu_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_cmp_ctl_wmr_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_async_por_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_peu_por_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_dmu_peu_wmr_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_l2_por_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_l2_wmr_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_niu_mac_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_niu_wmr_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_rst_por_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_rst_pwron_rst_sys2_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.rst_rst_wmr_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.state_ff.d0_0.d;
release tb_top.cpu.rst.rst_fsm_ctl.tr_flush_stop_ack_sys_ff.d0_0.d;
release tb_top.cpu.rst.rst_io_ctl.ccu_rst_change_io_ff.d0_0.d;
release tb_top.cpu.rst.rst_io_ctl.rst_rst_por_io_ff.d0_0.d;
release tb_top.cpu.rst.rst_io_ctl.rst_rst_pwron_rst_l_io_ff.d0_0.d;
release tb_top.cpu.rst.rst_io_ctl.rst_rst_wmr_io_ff.d0_0.d;
release tb_top.cpu.sii.clkgen_cmp.xcluster_header.alatch.d;
release tb_top.cpu.sii.clkgen_cmp.xcluster_header.blatch_divr.d;
release tb_top.cpu.sii.clkgen_cmp.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.sii.clkgen_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.sii.clkgen_cmp.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.sii.clkgen_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.sii.clkgen_io.xcluster_header.control_sig_sync.slow_cmp_sync_en_syncff.din_stg1.d;
release tb_top.cpu.sii.ilc0.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc0.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc0.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ilc1.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc1.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc1.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ilc2.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc2.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc2.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ilc3.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc3.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc3.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ilc4.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc4.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc4.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ilc5.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc5.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc5.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ilc6.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc6.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc6.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ilc7.reg_ilc_ild_addr_h.d0_0.d;
release tb_top.cpu.sii.ilc7.reg_ilc_ild_addr_lo.d0_0.d;
release tb_top.cpu.sii.ilc7.reg_ilc_ildq_rd_en.d0_0.d;
release tb_top.cpu.sii.ild0.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild0.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ild1.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild1.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ild2.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild2.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ild3.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild3.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ild4.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild4.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ild5.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild5.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ild6.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild6.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ild7.ff_sii_mb0_ild_fail.d0_0.d;
release tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_r.d0_0.d;
release tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_rr.d0_0.d;
release tb_top.cpu.sii.ild7.ff_sii_mb0_wdata_rrr.d0_0.d;
release tb_top.cpu.sii.ildq0.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq0.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq1.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq1.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq2.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq2.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq3.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq3.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq4.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq4.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq5.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq5.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq6.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq6.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq7.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ildq7.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.inc.reg_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.sii.inc.reg_mbist1_data_r.d0_0.d;
release tb_top.cpu.sii.inc.reg_mbist1_data_rr.d0_0.d;
release tb_top.cpu.sii.inc.reg_sii_mb0_ind_fail.d0_0.d;
release tb_top.cpu.sii.inc.reg_sii_mb0_wdata.d0_0.d;
release tb_top.cpu.sii.indq.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.indq.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipcc.reg_arb1.d0_0.d;
release tb_top.cpu.sii.ipcc.reg_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.sii.ipcc.reg_ncu_sii_ba01.d0_0.d;
release tb_top.cpu.sii.ipcc.reg_ncu_sii_ba23.d0_0.d;
release tb_top.cpu.sii.ipcc.reg_ncu_sii_ba45.d0_0.d;
release tb_top.cpu.sii.ipcc.reg_ncu_sii_ba67.d0_0.d;
release tb_top.cpu.sii.ipcc_dp.ff_mb0_wdata.d0_0.d;
release tb_top.cpu.sii.ipdbdq0_h.dff_din_hi.d0_0.d;
release tb_top.cpu.sii.ipdbdq0_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbdq0_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbdq0_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbdq0_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbdq1_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbdq1_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbdq1_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbdq1_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbhq0.dff_din_hi.d0_0.d;
release tb_top.cpu.sii.ipdbhq0.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbhq0.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbhq1.dff_din_hi.d0_0.d;
release tb_top.cpu.sii.ipdbhq1.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdbhq1.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq0_h.dff_din_hi.d0_0.d;
release tb_top.cpu.sii.ipdodq0_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq0_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq0_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq0_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq1_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq1_h.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq1_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdodq1_l.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdohq0.dff_din_hi.d0_0.d;
release tb_top.cpu.sii.ipdohq0.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdohq0.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdohq1.dff_din_hi.d0_0.d;
release tb_top.cpu.sii.ipdohq1.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.ipdohq1.dff_rd_en.d0_0.d;
release tb_top.cpu.sii.mb0.ild0_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ild1_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ild2_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ild3_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ild4_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ild5_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ild6_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ild7_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.ind_fail_reg.d0_0.d;
release tb_top.cpu.sii.mb0.wdata_reg.d0_0.d;
release tb_top.cpu.sii.mb1.data_pipe_reg1.d0_0.d;
release tb_top.cpu.sii.mb1.data_pipe_reg2.d0_0.d;
release tb_top.cpu.sii.mb1.data_pipe_reg3.d0_0.d;
release tb_top.cpu.sii.mb1.data_pipe_reg4.d0_0.d;
release tb_top.cpu.sii.mb1.data_pipe_reg5.d0_0.d;
release tb_top.cpu.sii.mb1.sel_pipe_reg1.d0_0.d;
release tb_top.cpu.sii.mb1.sel_pipe_reg2.d0_0.d;
release tb_top.cpu.sii.mb1.sel_reg.d0_0.d;
release tb_top.cpu.sii.mb1.wdata_reg.d0_0.d;
release tb_top.cpu.sii.mb1.wdata_reg2.d0_0.d;
release tb_top.cpu.sio.clkgen_cmp.xcluster_header.alatch.d;
release tb_top.cpu.sio.clkgen_cmp.xcluster_header.blatch_divr.d;
release tb_top.cpu.sio.clkgen_cmp.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.sio.clkgen_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.sio.clkgen_cmp.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.sio.clkgen_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.sio.clkgen_io.xcluster_header.control_sig_sync.slow_cmp_sync_en_syncff.din_stg1.d;
release tb_top.cpu.sio.mb0.data_pipe_reg1.d0_0.d;
release tb_top.cpu.sio.mb0.data_pipe_reg2.d0_0.d;
release tb_top.cpu.sio.mb0.data_pipe_reg3.d0_0.d;
release tb_top.cpu.sio.mb0.data_pipe_reg4.d0_0.d;
release tb_top.cpu.sio.mb0.read_data_pipe_reg.d0_0.d;
release tb_top.cpu.sio.mb0.wdata_reg.d0_0.d;
release tb_top.cpu.sio.mb1.data_pipe_reg1.d0_0.d;
release tb_top.cpu.sio.mb1.data_pipe_reg2.d0_0.d;
release tb_top.cpu.sio.mb1.data_pipe_reg3.d0_0.d;
release tb_top.cpu.sio.mb1.opd_sel_reg1.d0_0.d;
release tb_top.cpu.sio.mb1.opd_sel_reg2.d0_0.d;
release tb_top.cpu.sio.mb1.opd_sel_reg4.d0_0.d;
release tb_top.cpu.sio.mb1.read_data_pipe_reg.d0_0.d;
release tb_top.cpu.sio.mb1.sel_reg.d0_0.d;
release tb_top.cpu.sio.mb1.wdata_reg.d0_0.d;
release tb_top.cpu.sio.olddq00.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq01.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq10.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq11.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq20.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq21.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq30.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq31.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq40.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq41.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq50.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq51.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq60.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq61.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq70.dff_dout.d0_0.d;
release tb_top.cpu.sio.olddq71.dff_dout.d0_0.d;
release tb_top.cpu.sio.opcc.reg_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.sio.opcs0.reg_opdhqx_ue_bit.d0_0.d;
release tb_top.cpu.sio.opcs1.reg_opdhqx_ue_bit.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank01_data_opc1_h.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank01_data_opc1_l.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank23_data_opc1_h.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank23_data_opc1_l.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank45_data_opc1_h.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank45_data_opc1_l.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank67_data_opc1_h.d0_0.d;
release tb_top.cpu.sio.opdc.dff_bank67_data_opc1_l.d0_0.d;
release tb_top.cpu.sio.opdc.dff_mbist0145_data_h.d0_0.d;
release tb_top.cpu.sio.opdc.dff_mbist0145_data_l.d0_0.d;
release tb_top.cpu.sio.opdc.dff_mbist2367_data_h.d0_0.d;
release tb_top.cpu.sio.opdc.dff_mbist2367_data_l.d0_0.d;
release tb_top.cpu.sio.opddq00.dff_din_hi.d0_0.d;
release tb_top.cpu.sio.opddq00.dff_din_lo.d0_0.d;
release tb_top.cpu.sio.opddq00.dff_dout.d0_0.d;
release tb_top.cpu.sio.opddq01.dff_din_hi.d0_0.d;
release tb_top.cpu.sio.opddq01.dff_din_lo.d0_0.d;
release tb_top.cpu.sio.opddq01.dff_dout.d0_0.d;
release tb_top.cpu.sio.opddq10.dff_din_hi.d0_0.d;
release tb_top.cpu.sio.opddq10.dff_din_lo.d0_0.d;
release tb_top.cpu.sio.opddq10.dff_dout.d0_0.d;
release tb_top.cpu.sio.opddq11.dff_din_hi.d0_0.d;
release tb_top.cpu.sio.opddq11.dff_din_lo.d0_0.d;
release tb_top.cpu.sio.opddq11.dff_dout.d0_0.d;
release tb_top.cpu.sio.opdhq0.dff_din_hi.d0_0.d;
release tb_top.cpu.sio.opdhq0.dff_din_lo.d0_0.d;
release tb_top.cpu.sio.opdhq1.dff_din_hi.d0_0.d;
release tb_top.cpu.sio.opdhq1.dff_din_lo.d0_0.d;
release tb_top.cpu.sio.opds0.ff_opdhqxout.d0_0.d;
release tb_top.cpu.sio.opds0.ff_packet_data0_h.d0_0.d;
release tb_top.cpu.sio.opds0.ff_packet_data0_l.d0_0.d;
release tb_top.cpu.sio.opds0.ff_packet_data1_h.d0_0.d;
release tb_top.cpu.sio.opds0.ff_packet_data1_l.d0_0.d;
release tb_top.cpu.sio.opds1.ff_opdhqxout.d0_0.d;
release tb_top.cpu.sio.opds1.ff_packet_data0_h.d0_0.d;
release tb_top.cpu.sio.opds1.ff_packet_data0_l.d0_0.d;
release tb_top.cpu.sio.opds1.ff_packet_data1_h.d0_0.d;
release tb_top.cpu.sio.opds1.ff_packet_data1_l.d0_0.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.alatch.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.blatch_divr.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.spc0.clk_spc.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.spc0.dec.del.exu_clkenf.d0_0.d;
release tb_top.cpu.spc0.dec.del.fef.d0_0.d;
release tb_top.cpu.spc0.dec.del.pdisttidf.d0_0.d;
release tb_top.cpu.spc0.dec.del.tid_e.d0_0.d;
release tb_top.cpu.spc0.dec.del.tid_m.d0_0.d;
release tb_top.cpu.spc0.dec.del.truevalid_f.d0_0.d;
release tb_top.cpu.spc0.exu0.ect.fcce_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.ect.fgu_tid_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.ect.i_byp_lth.d0_0.d;
release tb_top.cpu.spc0.exu0.ect.i_estage_lth.d0_0.d;
release tb_top.cpu.spc0.exu0.ect.i_pwr0_lth.d0_0.d;
release tb_top.cpu.spc0.exu0.edp.i_asi0_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.edp.i_misc_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.irf.i_rd_control_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.irf.i_rd_control_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.irf.i_restore_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.irf.i_save_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.irf.i_wr_control_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.cansave_e2m2b2w.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.cleanwin_e2m2b2w.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.cwp_b2w.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.cwp_m2b.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.exception_report_m2b.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.i_rml_restore_en_ff.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.tid_p2d2e2m2b2w.d0_0.d;
release tb_top.cpu.spc0.exu0.rml.winblock_slot_tid_m2d2e2m.d0_0.d;
release tb_top.cpu.spc0.exu1.ect.fcce_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.ect.fgu_tid_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.ect.i_byp_lth.d0_0.d;
release tb_top.cpu.spc0.exu1.ect.i_estage_lth.d0_0.d;
release tb_top.cpu.spc0.exu1.ect.i_pwr0_lth.d0_0.d;
release tb_top.cpu.spc0.exu1.edp.i_asi0_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.edp.i_misc_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.irf.i_rd_control_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.irf.i_rd_control_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.irf.i_restore_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.irf.i_save_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.irf.i_wr_control_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.cansave_e2m2b2w.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.cleanwin_e2m2b2w.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.cwp_b2w.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.cwp_m2b.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.exception_report_m2b.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.i_rml_restore_en_ff.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.tid_p2d2e2m2b2w.d0_0.d;
release tb_top.cpu.spc0.exu1.rml.winblock_slot_tid_m2d2e2m.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.e_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.e_02.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fb_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fprs_frf_ctl.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fprs_rng.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fw_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fx1_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fx1_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fx2_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fx2_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fx3_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fx4_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.fx5_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.rng_6463.d0_0.d;
release tb_top.cpu.spc0.fgu.fac.rng_stg1.d0_0.d;
release tb_top.cpu.spc0.fgu.fad.e_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fad.e_01_extra.d0_0.d;
release tb_top.cpu.spc0.fgu.fdc.data_lth.d0_0.d;
release tb_top.cpu.spc0.fgu.fdc.ovlf_lth.d0_0.d;
release tb_top.cpu.spc0.fgu.fdc.xrnd_lth.d0_0.d;
release tb_top.cpu.spc0.fgu.fdd.ie_d00lthm1.d0_0.d;
release tb_top.cpu.spc0.fgu.fdd.ie_d00lthp1.d0_0.d;
release tb_top.cpu.spc0.fgu.fdd.ipte_clalth0.d0_0.d;
release tb_top.cpu.spc0.fgu.fdd.ipte_clalth1.d0_0.d;
release tb_top.cpu.spc0.fgu.fdd.isqe_cnt.d0_0.d;
release tb_top.cpu.spc0.fgu.fdd.isqe_flip.d0_0.d;
release tb_top.cpu.spc0.fgu.fgd.fx4_gsrtid.d0_0.d;
release tb_top.cpu.spc0.fgu.fic.fx2_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fb_05.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx1_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx2_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx2_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx2_02.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx2_05.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx3_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx3_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx3_02.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx3_03.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx3_05.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx3_06.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx4_00.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx4_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx4_02.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx5_01.d0_0.d;
release tb_top.cpu.spc0.fgu.fpc.fx5_02.d0_0.d;
release tb_top.cpu.spc0.fgu.fpe.fb_exp_res.d0_0.d;
release tb_top.cpu.spc0.fgu.fpe.fx1_fmtsel.d0_0.d;
release tb_top.cpu.spc0.fgu.fpe.fx2_aux.d0_0.d;
release tb_top.cpu.spc0.fgu.fpe.fx2_swp_sel.d0_0.d;
release tb_top.cpu.spc0.fgu.fpe.fx3_einty.d0_0.d;
release tb_top.cpu.spc0.fgu.fpe.fx4_einty.d0_0.d;
release tb_top.cpu.spc0.fgu.fpf.fb_nrd.d0_0.d;
release tb_top.cpu.spc0.fgu.fpf.fx2_fcc.d0_0.d;
release tb_top.cpu.spc0.fgu.fpf.fx3_fcc.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a0_be_ff.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a0_s_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a10_x_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a1_be_ff.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a1_s_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a2_be_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a2_s_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a32_x_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a3_be_ff.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a3_c_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a3_s_ff_a.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a4_c_hi_ff.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_a4_s_hi_ff.d0_0.d;
release tb_top.cpu.spc0.fgu.fpy.i_fx5_ff.d0_0.d;
release tb_top.cpu.spc0.fgu.frf.frf_read_ctl_in2ph2.d0_0.d;
release tb_top.cpu.spc0.fgu.frf.frf_write_input_ctl_in2fb.d0_0.d;
release tb_top.cpu.spc0.gkt.ipc.dff_ncu_pb.d0_0.d;
release tb_top.cpu.spc0.gkt.ipc.dff_pb_sel.d0_0.d;
release tb_top.cpu.spc0.gkt.ipc.dff_req_drop_latx.d0_0.d;
release tb_top.cpu.spc0.gkt.ipc.dff_unit_ndrop_pa.d0_0.d;
release tb_top.cpu.spc0.gkt.ipd.i_ifu_addr_v0_muxreg.d0_0.d;
release tb_top.cpu.spc0.gkt.ipd.i_mmu_addr_v0_muxreg.d0_0.d;
release tb_top.cpu.spc0.gkt.ipd.i_ncu_reg.d0_0.d;
release tb_top.cpu.spc0.gkt.ipd.i_req_li_reg.d0_0.d;
release tb_top.cpu.spc0.gkt.ipd.i_spu_addr_v0_muxreg.d0_0.d;
release tb_top.cpu.spc0.ifu_cmu.lsc.lsc_cpkt_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_cmu.lsd.paddr_lat.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.any_instr_v_c_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.br_misp_data_dup_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.br_misp_data_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.bus_first_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.ic_instr_v_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.inv_way1_bf_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.inv_way_bf_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_1_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_2_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.l2_cache_miss_in_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.mbist_output.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr0_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr1_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr2_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr3_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr4_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr5_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr6_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr7_pc_f_inc_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.thr_c_ic_disable_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.tid_dec_w_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_agc_ctl.wrway_bf_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_asi_ctl.rng_stg2_ctl.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_asi_ctl.rng_stg2_decctl.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_byp_dp.itb_data_for_cam.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_cms_ctl.rep_way_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.br_tid_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.itlb_probe_l_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.pstate_am_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_ftp_ctl.tid_dec_w_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.index_reg_i.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.quad_en_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.rdreq_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.way_c_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.way_f_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrreq_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_0_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_1_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_icd_cust.wrway_2_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.cache_way_hit_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tlb_cam_hit_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tte_tag_out_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.tte_u_bit_out_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_itc_ctl.itc_sel_demap_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_itc_ctl.tte1_lat.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_itd_dp.tte1_lat.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm0.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm1.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm2.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm3.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm4.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm5.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm6.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.ftu_tfc_ctl.tsm7.ignore_by_pass_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ftu.hdr.sram_header_instance.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq0.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq0.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq1.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq1.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq2.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq2.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq3.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq3.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq4.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq4.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq5.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq5.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq6.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq6.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq7.buff_clken_reg.d0_0.d;
release tb_top.cpu.spc0.ifu_ibu.ibq7.fetch_sig_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.ard.i_rngl_stg1_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.asc.ascl_vld_1.d0_0.d;
release tb_top.cpu.spc0.lsu.asc.hole_count.d0_0.d;
release tb_top.cpu.spc0.lsu.cic.dff_cpq_sel.d0_0.d;
release tb_top.cpu.spc0.lsu.dac.dff_baddr_b.d0_0.d;
release tb_top.cpu.spc0.lsu.dac.dff_endian_b.d0_0.d;
release tb_top.cpu.spc0.lsu.dac.dff_ld_sz_b.d0_0.d;
release tb_top.cpu.spc0.lsu.dca.dff_ctl_b.d0_0.d;
release tb_top.cpu.spc0.lsu.dca.dff_ctl_m_1.d0_0.d;
release tb_top.cpu.spc0.lsu.dca.lat_ctl_eb.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_asi_b.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_asi_m.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_excp_b.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_new_lru_w.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_pwr_mgmt.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_sba_par.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_tid_b.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_tid_e.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_tid_m.d0_0.d;
release tb_top.cpu.spc0.lsu.dcc.dff_tid_w.d0_0.d;
release tb_top.cpu.spc0.lsu.dcs.dff_context_m.d0_0.d;
release tb_top.cpu.spc0.lsu.dva.dff_din.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_inst_b.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_ld_inst_e.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_ld_lmq_en_b.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w2.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_ld_raw_w3.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_ld_sel.d0_0.d;
release tb_top.cpu.spc0.lsu.lmc.dff_thread_w.d0_0.d;
release tb_top.cpu.spc0.lsu.lru.dff_bit_en.d0_0.d;
release tb_top.cpu.spc0.lsu.lru.dff_din.d0_0.d;
release tb_top.cpu.spc0.lsu.pic.dff_asi_pm.d0_0.d;
release tb_top.cpu.spc0.lsu.pic.dff_asi_req.d0_0.d;
release tb_top.cpu.spc0.lsu.red.sram_header_instance.ff_io_cmp_sync_en.d0_0.d;
release tb_top.cpu.spc0.lsu.sbc.dff_cam_hit.d0_0.d;
release tb_top.cpu.spc0.lsu.sbc.dff_stb_err.d0_0.d;
release tb_top.cpu.spc0.lsu.sbc.dff_thread_b.d0_0.d;
release tb_top.cpu.spc0.lsu.sbc.dff_tid_m.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs0.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs1.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs2.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs3.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs4.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs5.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs6.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sbs7.dff_asi_pipe.d0_0.d;
release tb_top.cpu.spc0.lsu.sec.dff_cparity.d0_0.d;
release tb_top.cpu.spc0.lsu.sec.dff_st_sz.d0_0.d;
release tb_top.cpu.spc0.lsu.sed.dff_prty_bits.d0_0.d;
release tb_top.cpu.spc0.lsu.sed.dff_rd_data_0.d0_0.d;
release tb_top.cpu.spc0.lsu.sed.dff_rd_data_1.d0_0.d;
release tb_top.cpu.spc0.lsu.stb_cam.cam_tid_din.d0_0.d;
release tb_top.cpu.spc0.lsu.stb_cam.camwr_din.d0_0.d;
release tb_top.cpu.spc0.lsu.stb_cam.camwr_din.d0_0.d;
release tb_top.cpu.spc0.lsu.stb_ram.dff_din_lo.d0_0.d;
release tb_top.cpu.spc0.lsu.stb_ram.dff_wr_addr.d0_0.d;
release tb_top.cpu.spc0.lsu.tgd.dff_va_b.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.cache_way_hit_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.cam_ctl_lat.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.cam_ctl_lat.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.pa_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.page_size_mask_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.tlb_cam_hit_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.tte_data_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.tte_tag_out_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.tlb.tte_u_bit_out_reg.d0_0.d;
release tb_top.cpu.spc0.lsu.tlc.wr_vld_latch.d0_0.d;
release tb_top.cpu.spc0.lsu.tld.tte2_lat.d0_0.d;
release tb_top.cpu.spc0.mb0.cntl_reg.d0_0.d;
release tb_top.cpu.spc0.mb0.exp_stb_cam_hit_delay.d0_0.d;
release tb_top.cpu.spc0.mb0.input_signals_reg.d0_0.d;
release tb_top.cpu.spc0.mb0.pmen.d0_0.d;
release tb_top.cpu.spc0.mb1.cntl_reg.d0_0.d;
release tb_top.cpu.spc0.mb1.input_signals_reg.d0_0.d;
release tb_top.cpu.spc0.mb1.out_cmp_sel_reg.d0_0.d;
release tb_top.cpu.spc0.mb1.pmen.d0_0.d;
release tb_top.cpu.spc0.mb2.cntl_reg.d0_0.d;
release tb_top.cpu.spc0.mb2.input_signals_reg.d0_0.d;
release tb_top.cpu.spc0.mb2.pmen.d0_0.d;
release tb_top.cpu.spc0.mmu.ase.lsu_context_w_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.mbist_cmpsel_2_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.mbist_cmpsel_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.rd_tte_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.stg1_en_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.stg2_ctl_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.stg2_en_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.stg3_en_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.stg4_en_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.tag_access_tid_0_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.asi.tag_access_tid_1_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.gkt_hw0_lat0.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.hw4_stg_lat1.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.hw4_stg_lat2.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.m1_stg_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.m2_stg_lat2.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.m3_stg_lat1.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.rr_addr_hw2_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.htc.stg_hw3_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e0_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e1_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e2_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e3_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e4_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e5_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e6_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.e7_tte_reg_w40.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.reg_offsethw4_w27.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.reg_rangehw4_w55.d0_0.d;
release tb_top.cpu.spc0.mmu.htd.reg_tsbconf_m2_w39.d0_0.d;
release tb_top.cpu.spc0.mmu.mel0.ecc_lat.d0_0.d;
release tb_top.cpu.spc0.mmu.mel1.ecc_lat.d0_0.d;
release tb_top.cpu.spc0.msf0.bank2_lat.d0_0.d;
release tb_top.cpu.spc0.msf0.bank4_lat.d0_0.d;
release tb_top.cpu.spc0.pku.swl0.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl0.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl0.readyf.d0_0.d;
release tb_top.cpu.spc0.pku.swl1.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl1.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl1.readyf.d0_0.d;
release tb_top.cpu.spc0.pku.swl2.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl2.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl2.readyf.d0_0.d;
release tb_top.cpu.spc0.pku.swl3.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl3.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl3.readyf.d0_0.d;
release tb_top.cpu.spc0.pku.swl4.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl4.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl4.readyf.d0_0.d;
release tb_top.cpu.spc0.pku.swl5.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl5.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl5.readyf.d0_0.d;
release tb_top.cpu.spc0.pku.swl6.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl6.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl6.readyf.d0_0.d;
release tb_top.cpu.spc0.pku.swl7.not_annul_ds1_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl7.not_annul_ds2_f.d0_0.d;
release tb_top.cpu.spc0.pku.swl7.readyf.d0_0.d;
release tb_top.cpu.spc0.pmu.pmu_pct_ctl.asi.d0_0.d;
release tb_top.cpu.spc0.pmu.pmu_pct_ctl.events.d0_0.d;
release tb_top.cpu.spc0.pmu.pmu_pct_ctl.lsu_e2m.d0_0.d;
release tb_top.cpu.spc0.pmu.pmu_pct_ctl.lsutid.d0_0.d;
release tb_top.cpu.spc0.pmu.pmu_pct_ctl.pic_st.d0_0.d;
release tb_top.cpu.spc0.pmu.pmu_pct_ctl.pwrm.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.compare_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.mbist_cmpsel_2_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.mbist_cmpsel_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.rng_stg4.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.stg1_en_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.stg2_ctl_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.stg2_en_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.stg3_en_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.stg4_en_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.asi.wr_tid_dec_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.cep.asi_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls0.fast_tid_dec_b_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls0.hpriv_bar_or_ie_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls0.l1en_b2w_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls0.l_real_w_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls0.tid_b_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls0.tl_eq_0_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls1.fast_tid_dec_b_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls1.hpriv_bar_or_ie_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls1.l1en_b2w_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls1.l_real_w_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls1.tid_b_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.fls1.tl_eq_0_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.ras.s_dsfar_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.ras.tid0_b_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.ras.tid0_w1_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.ras.tid0_w_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.ras.tid1_b_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.ras.tid1_w1_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.ras.tid1_w_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.tca.dff_din_hi.d0_0.d;
release tb_top.cpu.spc0.tlu.tca.dff_rd_en.d0_0.d;
release tb_top.cpu.spc0.tlu.tca.dff_rd_en.d0_0.d;
release tb_top.cpu.spc0.tlu.tel0.ecc_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.tel1.ecc_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl0.gl_rest_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl0.l1en_per_thread_int_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl0.p_quiesce_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl0.pre_allow_don_ret_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl0.pre_allow_trap_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl0.stb_empty_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl0.tic_compare_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl1.gl_rest_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl1.l1en_per_thread_int_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl1.p_quiesce_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl1.pre_allow_don_ret_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl1.pre_allow_trap_lat.d0_0.d;
release tb_top.cpu.spc0.tlu.trl1.stb_empty_lat.d0_0.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.alatch.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.blatch_divr.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.ccu_div_ph_flop.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.tcu.clkgen_tcu_cmp.xcluster_header.observe_flops.obs_ff2.d;
release tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.clk_stopper.blatch.d;
release tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.por_syncff.din_stg1.d;
release tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.por_syncff.din_stg2.d;
release tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg1.d;
release tb_top.cpu.tcu.clkgen_tcu_io.xcluster_header.control_sig_sync.wmr_syncff.din_stg2.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_bnkstop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_cmpsync_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_l2tstop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_mcudrstop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_mcufbdstop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_mcuiostop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_mcustop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_soc0iostop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_soc0stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_soc1iostop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_soc2iostop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_soc3iostop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_soc3stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc0stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc1stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc2stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc3stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc4stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc5stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc6stop_reg.d0_0.d;
release tb_top.cpu.tcu.clkstp_ctl.clkstp_spc7stop_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.bank_avail_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.bank_enable_status_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.core_avail_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.core_enable_status_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.csr_mbist_mode_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.csr_ucb_data_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.dmo_ctl.dmo_dmodf_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.mbist_done_fail_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.mbist_done_reg.d0_0.d;
release tb_top.cpu.tcu.mbist_ctl.tcu_mbist_sync_en_reg.d0_0.d;
release tb_top.cpu.tcu.regs_ctl.spare_flops.d0_0.d;
release tb_top.cpu.tcu.regs_ctl.tcuregs_cmpiosync_reg.d0_0.d;
release tb_top.cpu.tcu.regs_ctl.tcuregs_ttstart_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk0_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk1_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk2_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk3_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk4_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk5_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk6_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopbnk7_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu0_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu1_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu2_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopmcu3_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc0_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc1_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc2_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopsoc3_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc0_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc1_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc2_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc3_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc4_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc5_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc6_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.clkseq_ctl.clkseq_stopspc7_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk0_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk1_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk1_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk2_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk2_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk3_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk4_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk4_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk5_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk5_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk6_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk6_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk7_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_bnk7_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t0_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t1_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t1_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t2_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t2_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t3_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t4_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t4_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t5_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t5_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t6_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t6_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t7_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_l2t7_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu0_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu1_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu1_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu2_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu2_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu3_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_mcu3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc0_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc1_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc2_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc3_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_soc3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc0_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc1_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc1_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc2_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc2_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc3_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc4_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc4_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc5_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc5_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc6_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc6_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc7_0.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_clk_stop_spc7_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu1_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu2_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_drclk_stop_mcu3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu1_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu2_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_mcu3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc0_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc1_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc2_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.sync_ff_ioclk_stop_soc3_1.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_cesq_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_cmpdrsync_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_cntdly_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_cntstart_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_cstopq48_nf_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_efcnt_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_efctl_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_enstat_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_flushclkstop_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_foffcnt_nf_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_fsreq_reg.d0_0.d;
release tb_top.cpu.tcu.sigmux_ctl.tcusig_rstsm_nf_reg.d0_0.d;

// 6260 signals released



// Reject list may follow...

// ccu path: instance=tb_top.cpu.ccu.ccu_core.align_pulse_cnt_bank5.U0.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.bf_sync1.xx0, model=cl_a1_msff_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.bf_sync1.xx1, model=cl_a1_msff_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.ccu_rst_sync_stable_ff.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.dr_sync_shift1.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.pll_div2_bnk6.U0, model=cl_a1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.pll_div2_bnk6.U1, model=cl_a1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.pll_div2_bnk6.U2, model=cl_a1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.pll_div3_bnk6.U0, model=cl_a1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.pll_div4_bnk6.U3, model=cl_a1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.rst_cnt_bank6.U1.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.rst_cnt_bank6.U2.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.rst_cnt_bank6.U4.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.rst_cnt_bank6.U5.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.sync2_shift.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_core.sys_cmp_sync_shift1.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_hm_wrapper.align_det.stg4.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_hm_wrapper.dr_reset_gen.dr_rst_n_ff.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_hm_wrapper.dr_reset_gen.pulse_wait.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.ccu_hm_wrapper.output_stg_eco2.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.clkgen_cmp.xcluster_header.alatch, model=cl_sc1_alatch_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.clkgen_cmp.xcluster_header.blatch_divr, model=cl_sc1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.clkgen_cmp.xcluster_header.ccu_div_ph_flop, model=cl_sc1_msff_1x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.clkgen_cmp.xcluster_header.clk_stopper.blatch, model=cl_sc1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.clkgen_cmp.xcluster_header.observe_flops.obs_ff2, model=cl_sc1_msff_1x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.clkgen_io.xcluster_header.clk_stopper.blatch, model=cl_sc1_blatch_4x, out=latout, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io2x_phase.clkout_tmp_0.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io2x_phase.flip_0.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io2x_phase.shift_bank_7.U1.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io2x_phase.shift_bank_7.U3.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io2x_phase.shift_bank_7.U5.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.cnt_bank5.U1.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.flip_0.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.phase_180_0.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.pre_phase_180_0.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.shift_bank_7.U1.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.shift_bank_7.U2.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.shift_bank_7.U5.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.gen_io_phase.shift_bank_7.U6.lib_inst, model=cl_a1_msff_arst_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.io_rstgen_blk.csr_ucb_rst_syncff.xx0, model=cl_a1_msff_4x, out=q, value=1
// ccu path: instance=tb_top.cpu.ccu.io_rstgen_blk.csr_ucb_rst_syncff.xx1, model=cl_a1_msff_4x, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.imaginary_vco_gen.pll_core, model=pll_core, out=vco_out, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x24, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x24, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x25, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x25, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x30, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x30, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x35, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x35, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x36, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x36, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x44, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.x8.x44, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.xd1.x24, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.xd1.x24, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.xd1.x43, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.xd1.x43, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.xd1.x44, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x1.xd1.x44, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x0.xb_0_, model=n2_core_pll_flop_reset2_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x0.xb_0_, model=n2_core_pll_flop_reset2_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x0.xb_1_, model=n2_core_pll_flop_reset2_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x0.xb_1_, model=n2_core_pll_flop_reset2_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x0.x17, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x0.x17, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x13, model=n2_core_pll_flop_reset2_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x13, model=n2_core_pll_flop_reset2_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x12, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x12, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x46, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x46, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x8, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x8, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x9, model=n2_core_pll_flop_reset2_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_0_.x2.x9, model=n2_core_pll_flop_reset2_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x13, model=n2_core_pll_flop_reset2_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x13, model=n2_core_pll_flop_reset2_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x12, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x12, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x22, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x22, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x45, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x45, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x46, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x46, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x8, model=n2_core_pll_flop_reset1_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x8, model=n2_core_pll_flop_reset1_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x9, model=n2_core_pll_flop_reset2_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x2_1_.x2.x9, model=n2_core_pll_flop_reset2_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x3.x0, model=n2_core_pll_flop_reset2_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x1.x3.x0, model=n2_core_pll_flop_reset2_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x0, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x0, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x19, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x19, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x20, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x20, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x23, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x23, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x3, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.x0.x3, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.xi72, model=n2_core_pll_flopderst_16x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.xi72, model=n2_core_pll_flopderst_16x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x2.xmxdel.x0.x0, model=decode, out=d, value=0001
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x0, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x0, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x19, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x19, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x20, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x20, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x23, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x23, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x3, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.x0.x3, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.xi72, model=n2_core_pll_flopderst_16x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.xi72, model=n2_core_pll_flopderst_16x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.x4.xmxdel.x0.x0, model=decode, out=d, value=0001
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.xd3.x24, model=n2_core_pll_tpm_gate2_cust, out=div_ck, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.xd3.x43, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.xd3.x43, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.xd3.x44, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.x6.xd3.x44, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x0, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x0, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x0, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x0, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x2, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x2, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x4, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x4, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x5, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x12.x5, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x0, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x0, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x2, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x2, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x4, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x4, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x5, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x15.x5, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x0, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x0, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x1, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x1, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x10, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x10, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x11, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x11, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x2, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x2, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x3, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x3, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x34, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x34, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x35, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x35, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x37, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x37, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x38, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x38, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x4, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x4, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x41, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x41, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x42, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x42, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x49, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x49, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x5, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x5, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x50, model=n2_core_pll_flop_reset_new_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x50, model=n2_core_pll_flop_reset_new_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x6, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x6, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x7, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x7, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x8, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x8, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x9, model=n2_core_pll_flop_reset_new_1x_cust, out=q, value=1
// invalid model: instance=tb_top.cpu.ccu.ccu_pll.xcharc.x16.x9, model=n2_core_pll_flop_reset_new_1x_cust, out=q_l, value=0
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x1.xccu_m0_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00111111111000111
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x1.xccu_m0_1, model=n2_clk_gl_cc_stage_4s4, out=stg5_out, value=1110
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x1.xccu_m0_2, model=n2_clk_gl_cc_stage_4s4, out=stg5_out, value=0001
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x11.xc1b_s4_0, model=n2_clk_gl_cc_stage_4s4, out=stg5_out, value=1011
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x12.xc1b_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000001111000
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x13.x35, model=n2_clk_gl_cc_stage_4s4, out=stg5_out, value=1111
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x14.xc2b_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000001111010
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x16.xc2t_s2_0, model=n2_clk_gl_cc_stage_8s2, out=stg5_out, value=00001101
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x19.xc2t_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000001101110
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x2.xc1t_s4_1, model=n2_clk_gl_cc_stage_4s4, out=stg5_out, value=0001
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x20.xc2t_s2_0, model=n2_clk_gl_cc_stage_8s2, out=stg5_out, value=00000001
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x21.xc2t_s2_0, model=n2_clk_gl_cc_stage_8s2, out=stg5_out, value=00001101
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x22.xc3t_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000001110000
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x24.xc2t_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000001111101
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x25.xc2t_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000000110101
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x26.xc3b_s1_2, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00010111000000000
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x27.xc2t_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000000000111
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x29.xc3b_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000110111000000
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x3.xc1t_s1_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000000001100000
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x5.xrst_m0_0, model=n2_clk_gl_cc_stage_17s1, out=stg1_out, value=00000001111111111
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x5.xrst_m0_1, model=n2_clk_gl_cc_stage_4s4, out=stg5_out, value=0011
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.x6.x6, model=n2_clk_gl_cc_stage_4s4, out=stg5_out, value=1101
// invalid model: instance=tb_top.cpu.n2_clk_gl_cust.n2_clk_gl_cc_stage_top_inst.xccu_align, model=n2_clk_gl_cc_stage_align, out=gclk_aligned, value=1
// invalid model: instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.i2cfdinteccchk11, model=ncu_eccchk11_ctl, out=co, value=11111
// invalid model: instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.i2cfdinteccchk11, model=ncu_eccchk11_ctl, out=dout, value=11111111111
// invalid model: instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.i2cfdioeccchk11, model=ncu_eccchk11_ctl, out=co, value=11111
// invalid model: instance=tb_top.cpu.ncu.ncu_fcd_ctl.ncu_i2cfcd_ctl.ncu_i2cfd_ctl.i2cfdioeccchk11, model=ncu_eccchk11_ctl, out=dout, value=11111111111
// invalid model: instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.c2ibufpioeccchk11, model=ncu_eccchk11_ctl, out=co, value=11111
// invalid model: instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.dmupio_ucb_buf.c2ibufpioeccchk11, model=ncu_eccchk11_ctl, out=dout, value=11111111111
// invalid model: instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_c2isd_ctl.c2isdeccchk6, model=ncu_eccchk6_ctl, out=co, value=11111
// invalid model: instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_c2isd_ctl.c2isdeccchk6, model=ncu_eccchk6_ctl, out=dout, value=111111
// invalid model: instance=tb_top.cpu.ncu.ncu_scd_ctl.ncu_c2iscd_ctl.ncu_c2isd_ctl.c2isdeccchk6, model=ncu_eccchk6_ctl, out=ue, value=1
// invalid model: instance=tb_top.cpu.spc0.ifu_ftu.ftu_itb_cust.array.cam, model=n2_tlb_tl_64x59_cam, out=tlb_cam_hit, value=1
// invalid model: instance=tb_top.cpu.spc0.lsu.tlb.array.cam, model=n2_tlb_tl_128x59_cam, out=tlb_cam_hit, value=1
// tisram_blb latout_l name: instance=tb_top.cpu.l2d0.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d0.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d1.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d1.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d2.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d2.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d3.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d3.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d4.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d4.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d5.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d5.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d6.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d6.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d7.ctr.tstmod.blb_read_c3_0.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2d7.ctr.tstmod.blb_read_c3_1.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t0.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t1.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t2.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t3.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t4.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t5.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t6.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad0.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad1.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad2.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank0.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank0.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank0.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank0.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank0.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank0.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank1.lat_reg_d_lft.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank1.lat_reg_d_rgt.d0_0, model=tisram_blb, out=latout_l, value=00000
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank1.lat_reg_en_lft.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank1.lat_reg_en_rgt.d0_0, model=tisram_blb, out=latout_l, value=00
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank1.lat_rid_lft.d0_0, model=tisram_blb, out=latout_l, value=0
// tisram_blb latout_l name: instance=tb_top.cpu.l2t7.tag.quad3.bank1.lat_rid_rgt.d0_0, model=tisram_blb, out=latout_l, value=0
// vcs barf: instance=tb_top.cpu.l2t0.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// vcs barf: instance=tb_top.cpu.l2t1.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// vcs barf: instance=tb_top.cpu.l2t2.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// vcs barf: instance=tb_top.cpu.l2t3.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// vcs barf: instance=tb_top.cpu.l2t4.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// vcs barf: instance=tb_top.cpu.l2t5.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// vcs barf: instance=tb_top.cpu.l2t6.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// vcs barf: instance=tb_top.cpu.l2t7.oque.ff_mux2_sel_c8_2.d0_0, model=dff, out=q, value=11111111111111111111111111111111111111
// x: instance=tb_top.cpu.ccu.csr_blk.rng_data_syncff.xx0, model=cl_a1_msff_4x, out=q, value=x
// x: instance=tb_top.cpu.ccu.csr_blk.rng_data_syncff.xx1, model=cl_a1_msff_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxn27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bsrxp27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.bscan.bstx19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd0.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu0.fbd1.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxn27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bsrxp27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.bscan.bstx19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd0.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu1.fbd1.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxn27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bsrxp27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.bscan.bstx19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd0.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu2.fbd1.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxn27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp20, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp21, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp22, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp23, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp24, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp25, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp26, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bsrxp27, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx00, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx01, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx02, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx03, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx04, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx05, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx06, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx07, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx08, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx09, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx10, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx11, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx12, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx13, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx14, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx15, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx16, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx17, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx18, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.bscan.bstx19, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd0.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf0.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf1.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf10.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf11.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf12.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf13.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf2.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf3.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf4.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf5.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf6.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf7.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf8.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat0, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat1, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat10, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat11, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat2, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat3, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat4, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat5, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat6, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat7, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat8, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mcu3.fbd1.frdbuf9.alat9, model=cl_dp1_alatch_4x, out=q, value=x
// x: instance=tb_top.cpu.mio.cell_17.ff_out, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mio.cell_2.ff_out, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mio.cell_209.ff_out, model=cl_sc1_bs_cell2_4x, out=q, value=x
// x: instance=tb_top.cpu.mio.muxsel.ff_1.d0_0, model=cl_sc1_msff_4x, out=q, value=x
// x: instance=tb_top.cpu.ncu.ncu_ssitop_ctl.ncu_ssisif_ctl.u_dff_io_jbi_ssi_miso_ff.d0_0, model=dff, out=q, value=x
// x: instance=tb_top.cpu.sii.ipcc.reg_dma_wr.d0_0, model=dff, out=q, value=x
// x: instance=tb_top.cpu.sii.ipcc_dp.ff_curhdri.d0_0, model=msffi_dp, out=q_l, value=xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx
// x: instance=tb_top.cpu.spc0.lsu.stb_cam.dff_out_addr.d0_0, model=dff, out=q, value=xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx
// x: instance=tb_top.cpu.spc0.lsu.stb_cam.dff_out_mask.d0_0, model=dff, out=q, value=xxxxxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_clkseqstat_reg.d0_0, model=dff, out=q, value=xx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_fusecoladdr_shift_reg.d0_0, model=dff, out=q, value=xxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_fusemode_shift_reg.d0_0, model=dff, out=q, value=xxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_fuserowaddr_shift_reg.d0_0, model=dff, out=q, value=xxxxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_idcode_reg.d0_0, model=dff, out=q, value=xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_lbist_bypass_shift_reg.d0_0, model=dff, out=q, value=xxxxxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_lbist_done_reg.d0_0, model=dff, out=q, value=xxxxxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_mbibypass_shift_reg.d0_0, model=dff, out=q, value=xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_mbist_get_done_fail_shift_reg.d0_0, model=dff, out=q, value=xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tap_mbist_result_reg.d0_0, model=dff, out=q, value=xx
// x: instance=tb_top.cpu.tcu.jtag_ctl.tcu_jtag_tap_ctl.bypass_ll_reg.d0_0, model=dff, out=q, value=x
// x: instance=tb_top.cpu.tcu.jtag_ctl.tcu_jtag_tap_ctl.bypass_reg.d0_0, model=dff, out=q, value=x
